library ieee;
use ieee.std_logic_1164.all;  

package koc_signal_pack is

    constant axi_resp_okay : std_logic_vector := "00";

end package;
