library ieee;
use ieee.std_logic_1164.all;

package main_pack is

	constant cpu_width : integer := 32;
	constant ram_size : integer := 1945;
	subtype word_type is std_logic_vector(cpu_width-1 downto 0);
	type ram_type is array(0 to ram_size-1) of word_type;
	function load_hex return ram_type;

end package;

package body main_pack is

	function load_hex return ram_type is
		variable ram_buffer : ram_type := (others=>(others=>'0'));
	begin
		ram_buffer(0) := X"3C1C1001";
		ram_buffer(1) := X"279C9E60";
		ram_buffer(2) := X"3C1D1000";
		ram_buffer(3) := X"27BD1E98";
		ram_buffer(4) := X"0C00012D";
		ram_buffer(5) := X"00000000";
		ram_buffer(6) := X"00000000";
		ram_buffer(7) := X"00000000";
		ram_buffer(8) := X"00000000";
		ram_buffer(9) := X"00000000";
		ram_buffer(10) := X"00000000";
		ram_buffer(11) := X"00000000";
		ram_buffer(12) := X"00000000";
		ram_buffer(13) := X"00000000";
		ram_buffer(14) := X"00000000";
		ram_buffer(15) := X"23BDFF98";
		ram_buffer(16) := X"AFA10010";
		ram_buffer(17) := X"AFA20014";
		ram_buffer(18) := X"AFA30018";
		ram_buffer(19) := X"AFA4001C";
		ram_buffer(20) := X"AFA50020";
		ram_buffer(21) := X"AFA60024";
		ram_buffer(22) := X"AFA70028";
		ram_buffer(23) := X"AFA8002C";
		ram_buffer(24) := X"AFA90030";
		ram_buffer(25) := X"AFAA0034";
		ram_buffer(26) := X"AFAB0038";
		ram_buffer(27) := X"AFAC003C";
		ram_buffer(28) := X"AFAD0040";
		ram_buffer(29) := X"AFAE0044";
		ram_buffer(30) := X"AFAF0048";
		ram_buffer(31) := X"AFB8004C";
		ram_buffer(32) := X"AFB90050";
		ram_buffer(33) := X"AFBF0054";
		ram_buffer(34) := X"401A7000";
		ram_buffer(35) := X"235AFFFC";
		ram_buffer(36) := X"AFBA0058";
		ram_buffer(37) := X"0000D810";
		ram_buffer(38) := X"AFBB005C";
		ram_buffer(39) := X"0000D812";
		ram_buffer(40) := X"AFBB0060";
		ram_buffer(41) := X"0C000103";
		ram_buffer(42) := X"23A50000";
		ram_buffer(43) := X"8FA10010";
		ram_buffer(44) := X"8FA20014";
		ram_buffer(45) := X"8FA30018";
		ram_buffer(46) := X"8FA4001C";
		ram_buffer(47) := X"8FA50020";
		ram_buffer(48) := X"8FA60024";
		ram_buffer(49) := X"8FA70028";
		ram_buffer(50) := X"8FA8002C";
		ram_buffer(51) := X"8FA90030";
		ram_buffer(52) := X"8FAA0034";
		ram_buffer(53) := X"8FAB0038";
		ram_buffer(54) := X"8FAC003C";
		ram_buffer(55) := X"8FAD0040";
		ram_buffer(56) := X"8FAE0044";
		ram_buffer(57) := X"8FAF0048";
		ram_buffer(58) := X"8FB8004C";
		ram_buffer(59) := X"8FB90050";
		ram_buffer(60) := X"8FBF0054";
		ram_buffer(61) := X"8FBA0058";
		ram_buffer(62) := X"8FBB005C";
		ram_buffer(63) := X"03600011";
		ram_buffer(64) := X"8FBB0060";
		ram_buffer(65) := X"03600013";
		ram_buffer(66) := X"23BD0068";
		ram_buffer(67) := X"341B0001";
		ram_buffer(68) := X"03400008";
		ram_buffer(69) := X"409B6000";
		ram_buffer(70) := X"40026000";
		ram_buffer(71) := X"03E00008";
		ram_buffer(72) := X"40846000";
		ram_buffer(73) := X"3C051000";
		ram_buffer(74) := X"24A50150";
		ram_buffer(75) := X"8CA60000";
		ram_buffer(76) := X"AC06003C";
		ram_buffer(77) := X"8CA60004";
		ram_buffer(78) := X"AC060040";
		ram_buffer(79) := X"8CA60008";
		ram_buffer(80) := X"AC060044";
		ram_buffer(81) := X"8CA6000C";
		ram_buffer(82) := X"03E00008";
		ram_buffer(83) := X"AC060048";
		ram_buffer(84) := X"3C1A1000";
		ram_buffer(85) := X"375A003C";
		ram_buffer(86) := X"03400008";
		ram_buffer(87) := X"00000000";
		ram_buffer(88) := X"00850019";
		ram_buffer(89) := X"00001012";
		ram_buffer(90) := X"00002010";
		ram_buffer(91) := X"03E00008";
		ram_buffer(92) := X"ACC40000";
		ram_buffer(93) := X"0000000C";
		ram_buffer(94) := X"03E00008";
		ram_buffer(95) := X"00000000";
		ram_buffer(96) := X"AC900000";
		ram_buffer(97) := X"AC910004";
		ram_buffer(98) := X"AC920008";
		ram_buffer(99) := X"AC93000C";
		ram_buffer(100) := X"AC940010";
		ram_buffer(101) := X"AC950014";
		ram_buffer(102) := X"AC960018";
		ram_buffer(103) := X"AC97001C";
		ram_buffer(104) := X"AC9E0020";
		ram_buffer(105) := X"AC9C0024";
		ram_buffer(106) := X"AC9D0028";
		ram_buffer(107) := X"AC9F002C";
		ram_buffer(108) := X"03E00008";
		ram_buffer(109) := X"34020000";
		ram_buffer(110) := X"8C900000";
		ram_buffer(111) := X"8C910004";
		ram_buffer(112) := X"8C920008";
		ram_buffer(113) := X"8C93000C";
		ram_buffer(114) := X"8C940010";
		ram_buffer(115) := X"8C950014";
		ram_buffer(116) := X"8C960018";
		ram_buffer(117) := X"8C97001C";
		ram_buffer(118) := X"8C9E0020";
		ram_buffer(119) := X"8C9C0024";
		ram_buffer(120) := X"8C9D0028";
		ram_buffer(121) := X"8C9F002C";
		ram_buffer(122) := X"03E00008";
		ram_buffer(123) := X"34A20000";
		ram_buffer(124) := X"27BDFFE0";
		ram_buffer(125) := X"AFBF001C";
		ram_buffer(126) := X"AFB10018";
		ram_buffer(127) := X"0C00061E";
		ram_buffer(128) := X"AFB00014";
		ram_buffer(129) := X"0C0006D0";
		ram_buffer(130) := X"24040001";
		ram_buffer(131) := X"3C021000";
		ram_buffer(132) := X"3C031000";
		ram_buffer(133) := X"24040005";
		ram_buffer(134) := X"AC601EB0";
		ram_buffer(135) := X"AC441EFC";
		ram_buffer(136) := X"8C441EFC";
		ram_buffer(137) := X"24631EB0";
		ram_buffer(138) := X"AC640004";
		ram_buffer(139) := X"8C640004";
		ram_buffer(140) := X"24421EFC";
		ram_buffer(141) := X"24840005";
		ram_buffer(142) := X"AC440004";
		ram_buffer(143) := X"8C450004";
		ram_buffer(144) := X"3C101000";
		ram_buffer(145) := X"3C111000";
		ram_buffer(146) := X"AC650008";
		ram_buffer(147) := X"26101D80";
		ram_buffer(148) := X"24030010";
		ram_buffer(149) := X"2631027C";
		ram_buffer(150) := X"2404000C";
		ram_buffer(151) := X"AC430008";
		ram_buffer(152) := X"0C00019D";
		ram_buffer(153) := X"AE110004";
		ram_buffer(154) := X"2404000C";
		ram_buffer(155) := X"0C00019D";
		ram_buffer(156) := X"AE110008";
		ram_buffer(157) := X"0C00009F";
		ram_buffer(158) := X"00000000";
		ram_buffer(159) := X"27BDFFC8";
		ram_buffer(160) := X"AFBF0034";
		ram_buffer(161) := X"AFB70030";
		ram_buffer(162) := X"AFB6002C";
		ram_buffer(163) := X"AFB50028";
		ram_buffer(164) := X"AFB40024";
		ram_buffer(165) := X"AFB30020";
		ram_buffer(166) := X"AFB2001C";
		ram_buffer(167) := X"AFB10018";
		ram_buffer(168) := X"AFB00014";
		ram_buffer(169) := X"3C02F000";
		ram_buffer(170) := X"8C420004";
		ram_buffer(171) := X"3C031000";
		ram_buffer(172) := X"3C041000";
		ram_buffer(173) := X"24841EFC";
		ram_buffer(174) := X"00021080";
		ram_buffer(175) := X"24631EB0";
		ram_buffer(176) := X"00431821";
		ram_buffer(177) := X"00441021";
		ram_buffer(178) := X"8C720000";
		ram_buffer(179) := X"8C550000";
		ram_buffer(180) := X"0C000655";
		ram_buffer(181) := X"3C141000";
		ram_buffer(182) := X"0C000709";
		ram_buffer(183) := X"0255882B";
		ram_buffer(184) := X"24500001";
		ram_buffer(185) := X"26941EBC";
		ram_buffer(186) := X"24160001";
		ram_buffer(187) := X"241701F3";
		ram_buffer(188) := X"0C0006FC";
		ram_buffer(189) := X"02002025";
		ram_buffer(190) := X"0C0006DE";
		ram_buffer(191) := X"26100001";
		ram_buffer(192) := X"0C0006D9";
		ram_buffer(193) := X"00000000";
		ram_buffer(194) := X"0C0006D4";
		ram_buffer(195) := X"00409825";
		ram_buffer(196) := X"12200019";
		ram_buffer(197) := X"02401825";
		ram_buffer(198) := X"10000009";
		ram_buffer(199) := X"00763004";
		ram_buffer(200) := X"8CA60000";
		ram_buffer(201) := X"00000000";
		ram_buffer(202) := X"24C60001";
		ram_buffer(203) := X"ACA60000";
		ram_buffer(204) := X"24630001";
		ram_buffer(205) := X"12A30010";
		ram_buffer(206) := X"00000000";
		ram_buffer(207) := X"00763004";
		ram_buffer(208) := X"00032880";
		ram_buffer(209) := X"02663824";
		ram_buffer(210) := X"10E0FFF9";
		ram_buffer(211) := X"02852821";
		ram_buffer(212) := X"8CA70000";
		ram_buffer(213) := X"00000000";
		ram_buffer(214) := X"14F7FFF1";
		ram_buffer(215) := X"00C23824";
		ram_buffer(216) := X"00062027";
		ram_buffer(217) := X"10E0000A";
		ram_buffer(218) := X"ACA00000";
		ram_buffer(219) := X"24630001";
		ram_buffer(220) := X"16A3FFF2";
		ram_buffer(221) := X"00441024";
		ram_buffer(222) := X"0C0006D0";
		ram_buffer(223) := X"00402025";
		ram_buffer(224) := X"0C0006EE";
		ram_buffer(225) := X"00000000";
		ram_buffer(226) := X"1000FFD9";
		ram_buffer(227) := X"00000000";
		ram_buffer(228) := X"1000FFE7";
		ram_buffer(229) := X"00461025";
		ram_buffer(230) := X"3C021000";
		ram_buffer(231) := X"3C031000";
		ram_buffer(232) := X"24040005";
		ram_buffer(233) := X"AC601EB0";
		ram_buffer(234) := X"AC441EFC";
		ram_buffer(235) := X"8C441EFC";
		ram_buffer(236) := X"24631EB0";
		ram_buffer(237) := X"AC640004";
		ram_buffer(238) := X"8C640004";
		ram_buffer(239) := X"24421EFC";
		ram_buffer(240) := X"24840005";
		ram_buffer(241) := X"AC440004";
		ram_buffer(242) := X"8C440004";
		ram_buffer(243) := X"00000000";
		ram_buffer(244) := X"AC640008";
		ram_buffer(245) := X"24030010";
		ram_buffer(246) := X"AC430008";
		ram_buffer(247) := X"03E00008";
		ram_buffer(248) := X"00000000";
		ram_buffer(249) := X"3C02F000";
		ram_buffer(250) := X"8C420004";
		ram_buffer(251) := X"3C031000";
		ram_buffer(252) := X"24631D8C";
		ram_buffer(253) := X"00021080";
		ram_buffer(254) := X"00431021";
		ram_buffer(255) := X"8C420000";
		ram_buffer(256) := X"24030002";
		ram_buffer(257) := X"03E00008";
		ram_buffer(258) := X"AC430000";
		ram_buffer(259) := X"27BDFFE0";
		ram_buffer(260) := X"AFBF001C";
		ram_buffer(261) := X"AFB20018";
		ram_buffer(262) := X"AFB10014";
		ram_buffer(263) := X"AFB00010";
		ram_buffer(264) := X"3C02F000";
		ram_buffer(265) := X"8C420004";
		ram_buffer(266) := X"00000000";
		ram_buffer(267) := X"00028100";
		ram_buffer(268) := X"02028021";
		ram_buffer(269) := X"00108080";
		ram_buffer(270) := X"26120004";
		ram_buffer(271) := X"3C111000";
		ram_buffer(272) := X"26311D98";
		ram_buffer(273) := X"02308021";
		ram_buffer(274) := X"8E020000";
		ram_buffer(275) := X"00000000";
		ram_buffer(276) := X"8C420004";
		ram_buffer(277) := X"00000000";
		ram_buffer(278) := X"2C430008";
		ram_buffer(279) := X"1060000F";
		ram_buffer(280) := X"00000000";
		ram_buffer(281) := X"000210C0";
		ram_buffer(282) := X"00521021";
		ram_buffer(283) := X"02221021";
		ram_buffer(284) := X"8C430000";
		ram_buffer(285) := X"8C440004";
		ram_buffer(286) := X"0060F809";
		ram_buffer(287) := X"00000000";
		ram_buffer(288) := X"8E020000";
		ram_buffer(289) := X"00000000";
		ram_buffer(290) := X"8C420004";
		ram_buffer(291) := X"00000000";
		ram_buffer(292) := X"2C430008";
		ram_buffer(293) := X"1460FFF3";
		ram_buffer(294) := X"00000000";
		ram_buffer(295) := X"8FBF001C";
		ram_buffer(296) := X"8FB20018";
		ram_buffer(297) := X"8FB10014";
		ram_buffer(298) := X"8FB00010";
		ram_buffer(299) := X"03E00008";
		ram_buffer(300) := X"27BD0020";
		ram_buffer(301) := X"27BDFFE0";
		ram_buffer(302) := X"AFBF001C";
		ram_buffer(303) := X"AFB20018";
		ram_buffer(304) := X"AFB10014";
		ram_buffer(305) := X"AFB00010";
		ram_buffer(306) := X"3C05F000";
		ram_buffer(307) := X"8CA20004";
		ram_buffer(308) := X"00000000";
		ram_buffer(309) := X"00021240";
		ram_buffer(310) := X"244301E8";
		ram_buffer(311) := X"3C021000";
		ram_buffer(312) := X"24421F08";
		ram_buffer(313) := X"00431021";
		ram_buffer(314) := X"0040E825";
		ram_buffer(315) := X"8CB00004";
		ram_buffer(316) := X"8CA60004";
		ram_buffer(317) := X"00000000";
		ram_buffer(318) := X"00062100";
		ram_buffer(319) := X"8CA50004";
		ram_buffer(320) := X"00861021";
		ram_buffer(321) := X"3C031000";
		ram_buffer(322) := X"3C071000";
		ram_buffer(323) := X"00021080";
		ram_buffer(324) := X"24631D98";
		ram_buffer(325) := X"24E71D8C";
		ram_buffer(326) := X"00052880";
		ram_buffer(327) := X"00624021";
		ram_buffer(328) := X"00A72821";
		ram_buffer(329) := X"24420004";
		ram_buffer(330) := X"3C09F002";
		ram_buffer(331) := X"00621021";
		ram_buffer(332) := X"ACA90000";
		ram_buffer(333) := X"25070044";
		ram_buffer(334) := X"3C05F001";
		ram_buffer(335) := X"AD050000";
		ram_buffer(336) := X"10470004";
		ram_buffer(337) := X"00402825";
		ram_buffer(338) := X"24A50008";
		ram_buffer(339) := X"14E5FFFE";
		ram_buffer(340) := X"ACA0FFF8";
		ram_buffer(341) := X"3C051000";
		ram_buffer(342) := X"24A503E4";
		ram_buffer(343) := X"AC450000";
		ram_buffer(344) := X"AC400004";
		ram_buffer(345) := X"00861021";
		ram_buffer(346) := X"00021080";
		ram_buffer(347) := X"00621821";
		ram_buffer(348) := X"8C620000";
		ram_buffer(349) := X"24030001";
		ram_buffer(350) := X"AC430000";
		ram_buffer(351) := X"1600000F";
		ram_buffer(352) := X"27838004";
		ram_buffer(353) := X"27828904";
		ram_buffer(354) := X"10620008";
		ram_buffer(355) := X"24660004";
		ram_buffer(356) := X"00463023";
		ram_buffer(357) := X"00063082";
		ram_buffer(358) := X"24C60001";
		ram_buffer(359) := X"00063080";
		ram_buffer(360) := X"00002825";
		ram_buffer(361) := X"0C000712";
		ram_buffer(362) := X"27848004";
		ram_buffer(363) := X"0C00007C";
		ram_buffer(364) := X"00000000";
		ram_buffer(365) := X"1000FFFF";
		ram_buffer(366) := X"00000000";
		ram_buffer(367) := X"0C00019D";
		ram_buffer(368) := X"2404000C";
		ram_buffer(369) := X"00101080";
		ram_buffer(370) := X"3C101000";
		ram_buffer(371) := X"26101D80";
		ram_buffer(372) := X"02028021";
		ram_buffer(373) := X"02008825";
		ram_buffer(374) := X"2412FFFF";
		ram_buffer(375) := X"24060004";
		ram_buffer(376) := X"02002825";
		ram_buffer(377) := X"0C000187";
		ram_buffer(378) := X"00002025";
		ram_buffer(379) := X"8E220000";
		ram_buffer(380) := X"00000000";
		ram_buffer(381) := X"1052FFFA";
		ram_buffer(382) := X"24060004";
		ram_buffer(383) := X"0C0001AD";
		ram_buffer(384) := X"00000000";
		ram_buffer(385) := X"8E220000";
		ram_buffer(386) := X"00000000";
		ram_buffer(387) := X"0040F809";
		ram_buffer(388) := X"00000000";
		ram_buffer(389) := X"1000FFE7";
		ram_buffer(390) := X"00000000";
		ram_buffer(391) := X"10C00013";
		ram_buffer(392) := X"00C51821";
		ram_buffer(393) := X"2406FFF0";
		ram_buffer(394) := X"00661024";
		ram_buffer(395) := X"0043182B";
		ram_buffer(396) := X"00031900";
		ram_buffer(397) := X"24420010";
		ram_buffer(398) := X"00A62824";
		ram_buffer(399) := X"00431821";
		ram_buffer(400) := X"40076000";
		ram_buffer(401) := X"40806000";
		ram_buffer(402) := X"10A30007";
		ram_buffer(403) := X"2484FF00";
		ram_buffer(404) := X"00A61024";
		ram_buffer(405) := X"AC820000";
		ram_buffer(406) := X"AC400000";
		ram_buffer(407) := X"24A50010";
		ram_buffer(408) := X"14A3FFFC";
		ram_buffer(409) := X"00A61024";
		ram_buffer(410) := X"40876000";
		ram_buffer(411) := X"03E00008";
		ram_buffer(412) := X"00000000";
		ram_buffer(413) := X"40066000";
		ram_buffer(414) := X"40806000";
		ram_buffer(415) := X"00001025";
		ram_buffer(416) := X"2483FF00";
		ram_buffer(417) := X"24050200";
		ram_buffer(418) := X"AC620000";
		ram_buffer(419) := X"AC400000";
		ram_buffer(420) := X"34440200";
		ram_buffer(421) := X"AC640000";
		ram_buffer(422) := X"AC800000";
		ram_buffer(423) := X"24420010";
		ram_buffer(424) := X"1445FFF9";
		ram_buffer(425) := X"00000000";
		ram_buffer(426) := X"40866000";
		ram_buffer(427) := X"03E00008";
		ram_buffer(428) := X"00000000";
		ram_buffer(429) := X"40066000";
		ram_buffer(430) := X"40806000";
		ram_buffer(431) := X"00000000";
		ram_buffer(432) := X"40076000";
		ram_buffer(433) := X"40806000";
		ram_buffer(434) := X"00001025";
		ram_buffer(435) := X"2403FF0C";
		ram_buffer(436) := X"24050200";
		ram_buffer(437) := X"AC620000";
		ram_buffer(438) := X"AC400000";
		ram_buffer(439) := X"34440200";
		ram_buffer(440) := X"AC640000";
		ram_buffer(441) := X"AC800000";
		ram_buffer(442) := X"24420010";
		ram_buffer(443) := X"1445FFF9";
		ram_buffer(444) := X"00000000";
		ram_buffer(445) := X"40876000";
		ram_buffer(446) := X"00000000";
		ram_buffer(447) := X"40076000";
		ram_buffer(448) := X"40806000";
		ram_buffer(449) := X"00001025";
		ram_buffer(450) := X"2403FF08";
		ram_buffer(451) := X"24050200";
		ram_buffer(452) := X"AC620000";
		ram_buffer(453) := X"AC400000";
		ram_buffer(454) := X"34440200";
		ram_buffer(455) := X"AC640000";
		ram_buffer(456) := X"AC800000";
		ram_buffer(457) := X"24420010";
		ram_buffer(458) := X"1445FFF9";
		ram_buffer(459) := X"00000000";
		ram_buffer(460) := X"40876000";
		ram_buffer(461) := X"00000000";
		ram_buffer(462) := X"40866000";
		ram_buffer(463) := X"03E00008";
		ram_buffer(464) := X"00000000";
		ram_buffer(465) := X"27BDFFB8";
		ram_buffer(466) := X"AFB60038";
		ram_buffer(467) := X"AFB50034";
		ram_buffer(468) := X"AFB40030";
		ram_buffer(469) := X"AFB20028";
		ram_buffer(470) := X"AFB10024";
		ram_buffer(471) := X"AFB00020";
		ram_buffer(472) := X"AFBF0044";
		ram_buffer(473) := X"AFBE0040";
		ram_buffer(474) := X"AFB7003C";
		ram_buffer(475) := X"AFB3002C";
		ram_buffer(476) := X"00809025";
		ram_buffer(477) := X"00A08825";
		ram_buffer(478) := X"00C08025";
		ram_buffer(479) := X"00E0A025";
		ram_buffer(480) := X"24150025";
		ram_buffer(481) := X"24160030";
		ram_buffer(482) := X"82050000";
		ram_buffer(483) := X"00000000";
		ram_buffer(484) := X"10A00009";
		ram_buffer(485) := X"00000000";
		ram_buffer(486) := X"10B50013";
		ram_buffer(487) := X"02402025";
		ram_buffer(488) := X"0220F809";
		ram_buffer(489) := X"26100001";
		ram_buffer(490) := X"82050000";
		ram_buffer(491) := X"00000000";
		ram_buffer(492) := X"14A0FFF9";
		ram_buffer(493) := X"00000000";
		ram_buffer(494) := X"8FBF0044";
		ram_buffer(495) := X"8FBE0040";
		ram_buffer(496) := X"8FB7003C";
		ram_buffer(497) := X"8FB60038";
		ram_buffer(498) := X"8FB50034";
		ram_buffer(499) := X"8FB40030";
		ram_buffer(500) := X"8FB3002C";
		ram_buffer(501) := X"8FB20028";
		ram_buffer(502) := X"8FB10024";
		ram_buffer(503) := X"8FB00020";
		ram_buffer(504) := X"03E00008";
		ram_buffer(505) := X"27BD0048";
		ram_buffer(506) := X"82040001";
		ram_buffer(507) := X"00000000";
		ram_buffer(508) := X"10960094";
		ram_buffer(509) := X"24060001";
		ram_buffer(510) := X"26100002";
		ram_buffer(511) := X"00003025";
		ram_buffer(512) := X"2482FFD0";
		ram_buffer(513) := X"304200FF";
		ram_buffer(514) := X"2C42000A";
		ram_buffer(515) := X"14400073";
		ram_buffer(516) := X"00001025";
		ram_buffer(517) := X"24030063";
		ram_buffer(518) := X"10830080";
		ram_buffer(519) := X"28830064";
		ram_buffer(520) := X"1460005F";
		ram_buffer(521) := X"24030073";
		ram_buffer(522) := X"108300C7";
		ram_buffer(523) := X"28830074";
		ram_buffer(524) := X"14600090";
		ram_buffer(525) := X"24030075";
		ram_buffer(526) := X"148300F0";
		ram_buffer(527) := X"24030078";
		ram_buffer(528) := X"8E840000";
		ram_buffer(529) := X"00000000";
		ram_buffer(530) := X"2C83000A";
		ram_buffer(531) := X"146001A7";
		ram_buffer(532) := X"26940004";
		ram_buffer(533) := X"24030001";
		ram_buffer(534) := X"00032880";
		ram_buffer(535) := X"00A31821";
		ram_buffer(536) := X"00031840";
		ram_buffer(537) := X"14600002";
		ram_buffer(538) := X"0083001B";
		ram_buffer(539) := X"0007000D";
		ram_buffer(540) := X"00002812";
		ram_buffer(541) := X"2CA5000A";
		ram_buffer(542) := X"10A0FFF8";
		ram_buffer(543) := X"00032880";
		ram_buffer(544) := X"1060001F";
		ram_buffer(545) := X"27AB0010";
		ram_buffer(546) := X"27A80010";
		ram_buffer(547) := X"00005025";
		ram_buffer(548) := X"240C000A";
		ram_buffer(549) := X"15800002";
		ram_buffer(550) := X"006C001B";
		ram_buffer(551) := X"0007000D";
		ram_buffer(552) := X"250B0001";
		ram_buffer(553) := X"24050057";
		ram_buffer(554) := X"00004812";
		ram_buffer(555) := X"00000000";
		ram_buffer(556) := X"00000000";
		ram_buffer(557) := X"14600002";
		ram_buffer(558) := X"0083001B";
		ram_buffer(559) := X"0007000D";
		ram_buffer(560) := X"00002010";
		ram_buffer(561) := X"00003812";
		ram_buffer(562) := X"15400003";
		ram_buffer(563) := X"01201825";
		ram_buffer(564) := X"18E0005F";
		ram_buffer(565) := X"00000000";
		ram_buffer(566) := X"28ED000A";
		ram_buffer(567) := X"11A00003";
		ram_buffer(568) := X"00A72821";
		ram_buffer(569) := X"24050030";
		ram_buffer(570) := X"00A72821";
		ram_buffer(571) := X"254A0001";
		ram_buffer(572) := X"11200003";
		ram_buffer(573) := X"A1050000";
		ram_buffer(574) := X"1000FFE6";
		ram_buffer(575) := X"01604025";
		ram_buffer(576) := X"14C0012D";
		ram_buffer(577) := X"A1600000";
		ram_buffer(578) := X"24170020";
		ram_buffer(579) := X"83B30010";
		ram_buffer(580) := X"00000000";
		ram_buffer(581) := X"1260017F";
		ram_buffer(582) := X"00000000";
		ram_buffer(583) := X"10400015";
		ram_buffer(584) := X"27A30011";
		ram_buffer(585) := X"10000004";
		ram_buffer(586) := X"24630001";
		ram_buffer(587) := X"10A00011";
		ram_buffer(588) := X"00A01025";
		ram_buffer(589) := X"24630001";
		ram_buffer(590) := X"8064FFFF";
		ram_buffer(591) := X"00000000";
		ram_buffer(592) := X"1480FFFA";
		ram_buffer(593) := X"2445FFFF";
		ram_buffer(594) := X"10A0000A";
		ram_buffer(595) := X"245EFFFE";
		ram_buffer(596) := X"02E02825";
		ram_buffer(597) := X"02402025";
		ram_buffer(598) := X"0220F809";
		ram_buffer(599) := X"27DEFFFF";
		ram_buffer(600) := X"27C20001";
		ram_buffer(601) := X"1C40FFFB";
		ram_buffer(602) := X"02E02825";
		ram_buffer(603) := X"1260FF86";
		ram_buffer(604) := X"00000000";
		ram_buffer(605) := X"27B70011";
		ram_buffer(606) := X"02602825";
		ram_buffer(607) := X"02402025";
		ram_buffer(608) := X"0220F809";
		ram_buffer(609) := X"26F70001";
		ram_buffer(610) := X"82F3FFFF";
		ram_buffer(611) := X"00000000";
		ram_buffer(612) := X"1660FFFA";
		ram_buffer(613) := X"02602825";
		ram_buffer(614) := X"1000FF7B";
		ram_buffer(615) := X"00000000";
		ram_buffer(616) := X"109500FE";
		ram_buffer(617) := X"24030058";
		ram_buffer(618) := X"10830096";
		ram_buffer(619) := X"00000000";
		ram_buffer(620) := X"1080FF81";
		ram_buffer(621) := X"00000000";
		ram_buffer(622) := X"1000FF73";
		ram_buffer(623) := X"00000000";
		ram_buffer(624) := X"2485FFD0";
		ram_buffer(625) := X"00021880";
		ram_buffer(626) := X"00621021";
		ram_buffer(627) := X"26100001";
		ram_buffer(628) := X"00021040";
		ram_buffer(629) := X"8204FFFF";
		ram_buffer(630) := X"00451021";
		ram_buffer(631) := X"308300FF";
		ram_buffer(632) := X"2465FFD0";
		ram_buffer(633) := X"2467FF9F";
		ram_buffer(634) := X"2CA5000A";
		ram_buffer(635) := X"14A0FFF4";
		ram_buffer(636) := X"2CE70006";
		ram_buffer(637) := X"2463FFBF";
		ram_buffer(638) := X"10E0000E";
		ram_buffer(639) := X"2C630006";
		ram_buffer(640) := X"2485FFA9";
		ram_buffer(641) := X"28A3000B";
		ram_buffer(642) := X"1460FFEF";
		ram_buffer(643) := X"00021880";
		ram_buffer(644) := X"24030063";
		ram_buffer(645) := X"1483FF82";
		ram_buffer(646) := X"28830064";
		ram_buffer(647) := X"82850003";
		ram_buffer(648) := X"02402025";
		ram_buffer(649) := X"0220F809";
		ram_buffer(650) := X"26940004";
		ram_buffer(651) := X"1000FF56";
		ram_buffer(652) := X"00000000";
		ram_buffer(653) := X"1060FF78";
		ram_buffer(654) := X"24030063";
		ram_buffer(655) := X"1000FFF1";
		ram_buffer(656) := X"2485FFC9";
		ram_buffer(657) := X"82040002";
		ram_buffer(658) := X"1000FF6D";
		ram_buffer(659) := X"26100003";
		ram_buffer(660) := X"152000D7";
		ram_buffer(661) := X"01005825";
		ram_buffer(662) := X"24E50030";
		ram_buffer(663) := X"250B0001";
		ram_buffer(664) := X"A1050000";
		ram_buffer(665) := X"10C0FFA8";
		ram_buffer(666) := X"A1600000";
		ram_buffer(667) := X"1000FFA7";
		ram_buffer(668) := X"24170030";
		ram_buffer(669) := X"24030064";
		ram_buffer(670) := X"1483FF43";
		ram_buffer(671) := X"00000000";
		ram_buffer(672) := X"8E850000";
		ram_buffer(673) := X"00000000";
		ram_buffer(674) := X"04A0010D";
		ram_buffer(675) := X"26940004";
		ram_buffer(676) := X"27A80010";
		ram_buffer(677) := X"28A3000A";
		ram_buffer(678) := X"14600110";
		ram_buffer(679) := X"00A03825";
		ram_buffer(680) := X"24030001";
		ram_buffer(681) := X"00032080";
		ram_buffer(682) := X"00831821";
		ram_buffer(683) := X"00031840";
		ram_buffer(684) := X"14600002";
		ram_buffer(685) := X"00A3001B";
		ram_buffer(686) := X"0007000D";
		ram_buffer(687) := X"00002012";
		ram_buffer(688) := X"2C84000A";
		ram_buffer(689) := X"1080FFF8";
		ram_buffer(690) := X"00032080";
		ram_buffer(691) := X"106000BE";
		ram_buffer(692) := X"01005825";
		ram_buffer(693) := X"00005025";
		ram_buffer(694) := X"240C000A";
		ram_buffer(695) := X"15800002";
		ram_buffer(696) := X"006C001B";
		ram_buffer(697) := X"0007000D";
		ram_buffer(698) := X"250B0001";
		ram_buffer(699) := X"24040057";
		ram_buffer(700) := X"00004812";
		ram_buffer(701) := X"00000000";
		ram_buffer(702) := X"00000000";
		ram_buffer(703) := X"14600002";
		ram_buffer(704) := X"00E3001B";
		ram_buffer(705) := X"0007000D";
		ram_buffer(706) := X"00003810";
		ram_buffer(707) := X"00002812";
		ram_buffer(708) := X"15400003";
		ram_buffer(709) := X"01201825";
		ram_buffer(710) := X"18A000D3";
		ram_buffer(711) := X"00000000";
		ram_buffer(712) := X"28AD000A";
		ram_buffer(713) := X"11A00003";
		ram_buffer(714) := X"00852021";
		ram_buffer(715) := X"24040030";
		ram_buffer(716) := X"00852021";
		ram_buffer(717) := X"254A0001";
		ram_buffer(718) := X"112000A3";
		ram_buffer(719) := X"A1040000";
		ram_buffer(720) := X"1000FFE6";
		ram_buffer(721) := X"01604025";
		ram_buffer(722) := X"8E970000";
		ram_buffer(723) := X"26940004";
		ram_buffer(724) := X"82E50000";
		ram_buffer(725) := X"00000000";
		ram_buffer(726) := X"10A000EA";
		ram_buffer(727) := X"26F30001";
		ram_buffer(728) := X"10400017";
		ram_buffer(729) := X"02601825";
		ram_buffer(730) := X"10000004";
		ram_buffer(731) := X"24630001";
		ram_buffer(732) := X"10C00013";
		ram_buffer(733) := X"00C01025";
		ram_buffer(734) := X"24630001";
		ram_buffer(735) := X"8064FFFF";
		ram_buffer(736) := X"00000000";
		ram_buffer(737) := X"1480FFFA";
		ram_buffer(738) := X"2446FFFF";
		ram_buffer(739) := X"10C0000C";
		ram_buffer(740) := X"245EFFFE";
		ram_buffer(741) := X"24050020";
		ram_buffer(742) := X"02402025";
		ram_buffer(743) := X"0220F809";
		ram_buffer(744) := X"27DEFFFF";
		ram_buffer(745) := X"27C20001";
		ram_buffer(746) := X"1C40FFFB";
		ram_buffer(747) := X"24050020";
		ram_buffer(748) := X"82E50000";
		ram_buffer(749) := X"00000000";
		ram_buffer(750) := X"10A0FEF3";
		ram_buffer(751) := X"00000000";
		ram_buffer(752) := X"02402025";
		ram_buffer(753) := X"0220F809";
		ram_buffer(754) := X"26730001";
		ram_buffer(755) := X"8265FFFF";
		ram_buffer(756) := X"00000000";
		ram_buffer(757) := X"10A0FEEC";
		ram_buffer(758) := X"02402025";
		ram_buffer(759) := X"0220F809";
		ram_buffer(760) := X"26730001";
		ram_buffer(761) := X"8265FFFF";
		ram_buffer(762) := X"00000000";
		ram_buffer(763) := X"14A0FFF5";
		ram_buffer(764) := X"02402025";
		ram_buffer(765) := X"1000FEE4";
		ram_buffer(766) := X"00000000";
		ram_buffer(767) := X"1483FEE2";
		ram_buffer(768) := X"00000000";
		ram_buffer(769) := X"8E850000";
		ram_buffer(770) := X"00000000";
		ram_buffer(771) := X"2CA30010";
		ram_buffer(772) := X"146000B4";
		ram_buffer(773) := X"26940004";
		ram_buffer(774) := X"24030001";
		ram_buffer(775) := X"00031900";
		ram_buffer(776) := X"14600002";
		ram_buffer(777) := X"00A3001B";
		ram_buffer(778) := X"0007000D";
		ram_buffer(779) := X"00003812";
		ram_buffer(780) := X"2CE70010";
		ram_buffer(781) := X"10E0FFF9";
		ram_buffer(782) := X"00000000";
		ram_buffer(783) := X"106000A5";
		ram_buffer(784) := X"00000000";
		ram_buffer(785) := X"24070058";
		ram_buffer(786) := X"27A90010";
		ram_buffer(787) := X"10870019";
		ram_buffer(788) := X"00005025";
		ram_buffer(789) := X"14600002";
		ram_buffer(790) := X"00A3001B";
		ram_buffer(791) := X"0007000D";
		ram_buffer(792) := X"00002810";
		ram_buffer(793) := X"00004012";
		ram_buffer(794) := X"15400003";
		ram_buffer(795) := X"00031902";
		ram_buffer(796) := X"19000082";
		ram_buffer(797) := X"00000000";
		ram_buffer(798) := X"290B000A";
		ram_buffer(799) := X"25240001";
		ram_buffer(800) := X"11600002";
		ram_buffer(801) := X"24070057";
		ram_buffer(802) := X"24070030";
		ram_buffer(803) := X"00E83821";
		ram_buffer(804) := X"254A0001";
		ram_buffer(805) := X"10600019";
		ram_buffer(806) := X"A1270000";
		ram_buffer(807) := X"1000FFED";
		ram_buffer(808) := X"00804825";
		ram_buffer(809) := X"10600078";
		ram_buffer(810) := X"25070030";
		ram_buffer(811) := X"01202025";
		ram_buffer(812) := X"00804825";
		ram_buffer(813) := X"14600002";
		ram_buffer(814) := X"00A3001B";
		ram_buffer(815) := X"0007000D";
		ram_buffer(816) := X"00002810";
		ram_buffer(817) := X"00004012";
		ram_buffer(818) := X"15400003";
		ram_buffer(819) := X"00031902";
		ram_buffer(820) := X"1900FFF4";
		ram_buffer(821) := X"00000000";
		ram_buffer(822) := X"290B000A";
		ram_buffer(823) := X"25240001";
		ram_buffer(824) := X"11600002";
		ram_buffer(825) := X"24070037";
		ram_buffer(826) := X"24070030";
		ram_buffer(827) := X"00E83821";
		ram_buffer(828) := X"254A0001";
		ram_buffer(829) := X"1460FFEE";
		ram_buffer(830) := X"A1270000";
		ram_buffer(831) := X"14C00030";
		ram_buffer(832) := X"A0800000";
		ram_buffer(833) := X"24170020";
		ram_buffer(834) := X"83B30010";
		ram_buffer(835) := X"00000000";
		ram_buffer(836) := X"12600084";
		ram_buffer(837) := X"00000000";
		ram_buffer(838) := X"10400015";
		ram_buffer(839) := X"27A30011";
		ram_buffer(840) := X"10000004";
		ram_buffer(841) := X"24630001";
		ram_buffer(842) := X"10A00011";
		ram_buffer(843) := X"00A01025";
		ram_buffer(844) := X"24630001";
		ram_buffer(845) := X"8064FFFF";
		ram_buffer(846) := X"00000000";
		ram_buffer(847) := X"1480FFFA";
		ram_buffer(848) := X"2445FFFF";
		ram_buffer(849) := X"10A0000A";
		ram_buffer(850) := X"245EFFFE";
		ram_buffer(851) := X"02E02825";
		ram_buffer(852) := X"02402025";
		ram_buffer(853) := X"0220F809";
		ram_buffer(854) := X"27DEFFFF";
		ram_buffer(855) := X"27C20001";
		ram_buffer(856) := X"1C40FFFB";
		ram_buffer(857) := X"02E02825";
		ram_buffer(858) := X"1260FE87";
		ram_buffer(859) := X"00000000";
		ram_buffer(860) := X"27B70011";
		ram_buffer(861) := X"02602825";
		ram_buffer(862) := X"02402025";
		ram_buffer(863) := X"0220F809";
		ram_buffer(864) := X"26F70001";
		ram_buffer(865) := X"82F3FFFF";
		ram_buffer(866) := X"00000000";
		ram_buffer(867) := X"1660FFFA";
		ram_buffer(868) := X"02602825";
		ram_buffer(869) := X"1000FE7C";
		ram_buffer(870) := X"00000000";
		ram_buffer(871) := X"24050025";
		ram_buffer(872) := X"0220F809";
		ram_buffer(873) := X"02402025";
		ram_buffer(874) := X"1000FE77";
		ram_buffer(875) := X"00000000";
		ram_buffer(876) := X"1000FEB8";
		ram_buffer(877) := X"01604025";
		ram_buffer(878) := X"1000FED4";
		ram_buffer(879) := X"24170030";
		ram_buffer(880) := X"1000FFD1";
		ram_buffer(881) := X"24170030";
		ram_buffer(882) := X"10C00039";
		ram_buffer(883) := X"A1600000";
		ram_buffer(884) := X"24170030";
		ram_buffer(885) := X"83B30010";
		ram_buffer(886) := X"00000000";
		ram_buffer(887) := X"12600045";
		ram_buffer(888) := X"00000000";
		ram_buffer(889) := X"10400015";
		ram_buffer(890) := X"27A30011";
		ram_buffer(891) := X"10000004";
		ram_buffer(892) := X"24630001";
		ram_buffer(893) := X"10A00011";
		ram_buffer(894) := X"00A01025";
		ram_buffer(895) := X"24630001";
		ram_buffer(896) := X"8064FFFF";
		ram_buffer(897) := X"00000000";
		ram_buffer(898) := X"1480FFFA";
		ram_buffer(899) := X"2445FFFF";
		ram_buffer(900) := X"10A0000A";
		ram_buffer(901) := X"245EFFFE";
		ram_buffer(902) := X"02E02825";
		ram_buffer(903) := X"02402025";
		ram_buffer(904) := X"0220F809";
		ram_buffer(905) := X"27DEFFFF";
		ram_buffer(906) := X"27C20001";
		ram_buffer(907) := X"1C40FFFB";
		ram_buffer(908) := X"02E02825";
		ram_buffer(909) := X"1260FE54";
		ram_buffer(910) := X"00000000";
		ram_buffer(911) := X"27B70011";
		ram_buffer(912) := X"02602825";
		ram_buffer(913) := X"02402025";
		ram_buffer(914) := X"0220F809";
		ram_buffer(915) := X"26F70001";
		ram_buffer(916) := X"82F3FFFF";
		ram_buffer(917) := X"00000000";
		ram_buffer(918) := X"1660FFFA";
		ram_buffer(919) := X"02602825";
		ram_buffer(920) := X"1000FE49";
		ram_buffer(921) := X"00000000";
		ram_buffer(922) := X"1120000D";
		ram_buffer(923) := X"24A40030";
		ram_buffer(924) := X"01005825";
		ram_buffer(925) := X"1000FF19";
		ram_buffer(926) := X"01604025";
		ram_buffer(927) := X"1460000E";
		ram_buffer(928) := X"01202025";
		ram_buffer(929) := X"25070030";
		ram_buffer(930) := X"25240001";
		ram_buffer(931) := X"A1270000";
		ram_buffer(932) := X"10C0FF9C";
		ram_buffer(933) := X"A0800000";
		ram_buffer(934) := X"1000FF9B";
		ram_buffer(935) := X"24170030";
		ram_buffer(936) := X"250B0001";
		ram_buffer(937) := X"A1040000";
		ram_buffer(938) := X"14C0FFC9";
		ram_buffer(939) := X"A1600000";
		ram_buffer(940) := X"1000FFC8";
		ram_buffer(941) := X"24170020";
		ram_buffer(942) := X"1000FF66";
		ram_buffer(943) := X"00804825";
		ram_buffer(944) := X"2403002D";
		ram_buffer(945) := X"00052823";
		ram_buffer(946) := X"A3A30010";
		ram_buffer(947) := X"1000FEF1";
		ram_buffer(948) := X"27A80011";
		ram_buffer(949) := X"1000FF89";
		ram_buffer(950) := X"27A40010";
		ram_buffer(951) := X"1000FEFD";
		ram_buffer(952) := X"24030001";
		ram_buffer(953) := X"1000FF57";
		ram_buffer(954) := X"24030001";
		ram_buffer(955) := X"1000FE66";
		ram_buffer(956) := X"24030001";
		ram_buffer(957) := X"1040FE24";
		ram_buffer(958) := X"245EFFFF";
		ram_buffer(959) := X"1000FFC7";
		ram_buffer(960) := X"02E02825";
		ram_buffer(961) := X"1040FE20";
		ram_buffer(962) := X"245EFFFF";
		ram_buffer(963) := X"1000FF22";
		ram_buffer(964) := X"24050020";
		ram_buffer(965) := X"1040FE1C";
		ram_buffer(966) := X"245EFFFF";
		ram_buffer(967) := X"1000FE8D";
		ram_buffer(968) := X"02E02825";
		ram_buffer(969) := X"1040FE18";
		ram_buffer(970) := X"245EFFFF";
		ram_buffer(971) := X"1000FF88";
		ram_buffer(972) := X"02E02825";
		ram_buffer(973) := X"AF858008";
		ram_buffer(974) := X"03E00008";
		ram_buffer(975) := X"AF848004";
		ram_buffer(976) := X"27BDFFE0";
		ram_buffer(977) := X"27A20024";
		ram_buffer(978) := X"AFA50024";
		ram_buffer(979) := X"AFA60028";
		ram_buffer(980) := X"8F858008";
		ram_buffer(981) := X"00803025";
		ram_buffer(982) := X"8F848004";
		ram_buffer(983) := X"AFA7002C";
		ram_buffer(984) := X"00403825";
		ram_buffer(985) := X"AFBF001C";
		ram_buffer(986) := X"0C0001D1";
		ram_buffer(987) := X"AFA20010";
		ram_buffer(988) := X"8FBF001C";
		ram_buffer(989) := X"00000000";
		ram_buffer(990) := X"03E00008";
		ram_buffer(991) := X"27BD0020";
		ram_buffer(992) := X"27BDFFC0";
		ram_buffer(993) := X"AFB50034";
		ram_buffer(994) := X"27B50048";
		ram_buffer(995) := X"AFB3002C";
		ram_buffer(996) := X"AFB20028";
		ram_buffer(997) := X"AFB10024";
		ram_buffer(998) := X"AFBF003C";
		ram_buffer(999) := X"AFB60038";
		ram_buffer(1000) := X"AFB40030";
		ram_buffer(1001) := X"AFB00020";
		ram_buffer(1002) := X"00801825";
		ram_buffer(1003) := X"00A08825";
		ram_buffer(1004) := X"AFA60048";
		ram_buffer(1005) := X"AFA7004C";
		ram_buffer(1006) := X"AFB5001C";
		ram_buffer(1007) := X"24120025";
		ram_buffer(1008) := X"24130030";
		ram_buffer(1009) := X"82220000";
		ram_buffer(1010) := X"00000000";
		ram_buffer(1011) := X"10400009";
		ram_buffer(1012) := X"00000000";
		ram_buffer(1013) := X"10520012";
		ram_buffer(1014) := X"00000000";
		ram_buffer(1015) := X"A0620000";
		ram_buffer(1016) := X"26310001";
		ram_buffer(1017) := X"82220000";
		ram_buffer(1018) := X"00000000";
		ram_buffer(1019) := X"1440FFF9";
		ram_buffer(1020) := X"24630001";
		ram_buffer(1021) := X"A0600000";
		ram_buffer(1022) := X"8FBF003C";
		ram_buffer(1023) := X"8FB60038";
		ram_buffer(1024) := X"8FB50034";
		ram_buffer(1025) := X"8FB40030";
		ram_buffer(1026) := X"8FB3002C";
		ram_buffer(1027) := X"8FB20028";
		ram_buffer(1028) := X"8FB10024";
		ram_buffer(1029) := X"8FB00020";
		ram_buffer(1030) := X"03E00008";
		ram_buffer(1031) := X"27BD0040";
		ram_buffer(1032) := X"82240001";
		ram_buffer(1033) := X"00000000";
		ram_buffer(1034) := X"10930090";
		ram_buffer(1035) := X"24070001";
		ram_buffer(1036) := X"26310002";
		ram_buffer(1037) := X"00003825";
		ram_buffer(1038) := X"2482FFD0";
		ram_buffer(1039) := X"304200FF";
		ram_buffer(1040) := X"2C42000A";
		ram_buffer(1041) := X"14400043";
		ram_buffer(1042) := X"00008025";
		ram_buffer(1043) := X"24020063";
		ram_buffer(1044) := X"10820050";
		ram_buffer(1045) := X"28820064";
		ram_buffer(1046) := X"1440007C";
		ram_buffer(1047) := X"24020073";
		ram_buffer(1048) := X"108200C3";
		ram_buffer(1049) := X"28820074";
		ram_buffer(1050) := X"1440008C";
		ram_buffer(1051) := X"24020075";
		ram_buffer(1052) := X"148200ED";
		ram_buffer(1053) := X"24020078";
		ram_buffer(1054) := X"8EA40000";
		ram_buffer(1055) := X"00000000";
		ram_buffer(1056) := X"2C82000A";
		ram_buffer(1057) := X"144001AA";
		ram_buffer(1058) := X"26B50004";
		ram_buffer(1059) := X"24020001";
		ram_buffer(1060) := X"00022880";
		ram_buffer(1061) := X"00A21021";
		ram_buffer(1062) := X"00021040";
		ram_buffer(1063) := X"14400002";
		ram_buffer(1064) := X"0082001B";
		ram_buffer(1065) := X"0007000D";
		ram_buffer(1066) := X"00002812";
		ram_buffer(1067) := X"2CA5000A";
		ram_buffer(1068) := X"10A0FFF8";
		ram_buffer(1069) := X"00022880";
		ram_buffer(1070) := X"1040003B";
		ram_buffer(1071) := X"27AB0010";
		ram_buffer(1072) := X"27A80010";
		ram_buffer(1073) := X"00005025";
		ram_buffer(1074) := X"240C000A";
		ram_buffer(1075) := X"15800002";
		ram_buffer(1076) := X"004C001B";
		ram_buffer(1077) := X"0007000D";
		ram_buffer(1078) := X"250B0001";
		ram_buffer(1079) := X"24050057";
		ram_buffer(1080) := X"00004812";
		ram_buffer(1081) := X"00000000";
		ram_buffer(1082) := X"00000000";
		ram_buffer(1083) := X"14400002";
		ram_buffer(1084) := X"0082001B";
		ram_buffer(1085) := X"0007000D";
		ram_buffer(1086) := X"00002010";
		ram_buffer(1087) := X"00003012";
		ram_buffer(1088) := X"15400003";
		ram_buffer(1089) := X"01201025";
		ram_buffer(1090) := X"18C0005B";
		ram_buffer(1091) := X"00000000";
		ram_buffer(1092) := X"28CD000A";
		ram_buffer(1093) := X"11A00003";
		ram_buffer(1094) := X"00A62821";
		ram_buffer(1095) := X"24050030";
		ram_buffer(1096) := X"00A62821";
		ram_buffer(1097) := X"254A0001";
		ram_buffer(1098) := X"1120001F";
		ram_buffer(1099) := X"A1050000";
		ram_buffer(1100) := X"1000FFE6";
		ram_buffer(1101) := X"01604025";
		ram_buffer(1102) := X"2485FFD0";
		ram_buffer(1103) := X"00101080";
		ram_buffer(1104) := X"00508021";
		ram_buffer(1105) := X"26310001";
		ram_buffer(1106) := X"00108040";
		ram_buffer(1107) := X"8224FFFF";
		ram_buffer(1108) := X"02058021";
		ram_buffer(1109) := X"308200FF";
		ram_buffer(1110) := X"2445FFD0";
		ram_buffer(1111) := X"2446FF9F";
		ram_buffer(1112) := X"2CA5000A";
		ram_buffer(1113) := X"14A0FFF4";
		ram_buffer(1114) := X"2CC60006";
		ram_buffer(1115) := X"2442FFBF";
		ram_buffer(1116) := X"10C00032";
		ram_buffer(1117) := X"2C420006";
		ram_buffer(1118) := X"2485FFA9";
		ram_buffer(1119) := X"28A2000B";
		ram_buffer(1120) := X"1440FFEF";
		ram_buffer(1121) := X"00101080";
		ram_buffer(1122) := X"24020063";
		ram_buffer(1123) := X"1482FFB2";
		ram_buffer(1124) := X"28820064";
		ram_buffer(1125) := X"8EA20000";
		ram_buffer(1126) := X"24630001";
		ram_buffer(1127) := X"A062FFFF";
		ram_buffer(1128) := X"1000FF88";
		ram_buffer(1129) := X"26B50004";
		ram_buffer(1130) := X"14E00109";
		ram_buffer(1131) := X"A1600000";
		ram_buffer(1132) := X"24050020";
		ram_buffer(1133) := X"83B40010";
		ram_buffer(1134) := X"00000000";
		ram_buffer(1135) := X"1280014A";
		ram_buffer(1136) := X"00000000";
		ram_buffer(1137) := X"12000013";
		ram_buffer(1138) := X"27A20011";
		ram_buffer(1139) := X"10000004";
		ram_buffer(1140) := X"24420001";
		ram_buffer(1141) := X"10C0000F";
		ram_buffer(1142) := X"00C08025";
		ram_buffer(1143) := X"24420001";
		ram_buffer(1144) := X"8044FFFF";
		ram_buffer(1145) := X"00000000";
		ram_buffer(1146) := X"1480FFFA";
		ram_buffer(1147) := X"2606FFFF";
		ram_buffer(1148) := X"10C00008";
		ram_buffer(1149) := X"2610FFFE";
		ram_buffer(1150) := X"06000145";
		ram_buffer(1151) := X"00000000";
		ram_buffer(1152) := X"26100001";
		ram_buffer(1153) := X"00602025";
		ram_buffer(1154) := X"0C000712";
		ram_buffer(1155) := X"02003025";
		ram_buffer(1156) := X"00501821";
		ram_buffer(1157) := X"27A20011";
		ram_buffer(1158) := X"24630001";
		ram_buffer(1159) := X"24420001";
		ram_buffer(1160) := X"A074FFFF";
		ram_buffer(1161) := X"8054FFFF";
		ram_buffer(1162) := X"00000000";
		ram_buffer(1163) := X"1680FFFB";
		ram_buffer(1164) := X"24630001";
		ram_buffer(1165) := X"1000FF63";
		ram_buffer(1166) := X"2463FFFF";
		ram_buffer(1167) := X"1040FF84";
		ram_buffer(1168) := X"24020063";
		ram_buffer(1169) := X"1000FFCD";
		ram_buffer(1170) := X"2485FFC9";
		ram_buffer(1171) := X"109200DB";
		ram_buffer(1172) := X"24020058";
		ram_buffer(1173) := X"10820076";
		ram_buffer(1174) := X"00000000";
		ram_buffer(1175) := X"1080FF65";
		ram_buffer(1176) := X"00000000";
		ram_buffer(1177) := X"1000FF57";
		ram_buffer(1178) := X"00000000";
		ram_buffer(1179) := X"82240002";
		ram_buffer(1180) := X"1000FF71";
		ram_buffer(1181) := X"26310003";
		ram_buffer(1182) := X"152000D3";
		ram_buffer(1183) := X"01005825";
		ram_buffer(1184) := X"24C50030";
		ram_buffer(1185) := X"250B0001";
		ram_buffer(1186) := X"A1050000";
		ram_buffer(1187) := X"10E0FFC8";
		ram_buffer(1188) := X"A1600000";
		ram_buffer(1189) := X"1000FFC7";
		ram_buffer(1190) := X"24050030";
		ram_buffer(1191) := X"24020064";
		ram_buffer(1192) := X"1482FF48";
		ram_buffer(1193) := X"00000000";
		ram_buffer(1194) := X"8EA50000";
		ram_buffer(1195) := X"00000000";
		ram_buffer(1196) := X"04A00106";
		ram_buffer(1197) := X"26B50004";
		ram_buffer(1198) := X"27A80010";
		ram_buffer(1199) := X"28A2000A";
		ram_buffer(1200) := X"14400117";
		ram_buffer(1201) := X"00A03025";
		ram_buffer(1202) := X"24020001";
		ram_buffer(1203) := X"00022080";
		ram_buffer(1204) := X"00821021";
		ram_buffer(1205) := X"00021040";
		ram_buffer(1206) := X"14400002";
		ram_buffer(1207) := X"00A2001B";
		ram_buffer(1208) := X"0007000D";
		ram_buffer(1209) := X"00002012";
		ram_buffer(1210) := X"2C84000A";
		ram_buffer(1211) := X"1080FFF8";
		ram_buffer(1212) := X"00022080";
		ram_buffer(1213) := X"104000BA";
		ram_buffer(1214) := X"01005825";
		ram_buffer(1215) := X"00005025";
		ram_buffer(1216) := X"240C000A";
		ram_buffer(1217) := X"15800002";
		ram_buffer(1218) := X"004C001B";
		ram_buffer(1219) := X"0007000D";
		ram_buffer(1220) := X"250B0001";
		ram_buffer(1221) := X"24040057";
		ram_buffer(1222) := X"00004812";
		ram_buffer(1223) := X"00000000";
		ram_buffer(1224) := X"00000000";
		ram_buffer(1225) := X"14400002";
		ram_buffer(1226) := X"00C2001B";
		ram_buffer(1227) := X"0007000D";
		ram_buffer(1228) := X"00003010";
		ram_buffer(1229) := X"00002812";
		ram_buffer(1230) := X"15400003";
		ram_buffer(1231) := X"01201025";
		ram_buffer(1232) := X"18A000CC";
		ram_buffer(1233) := X"00000000";
		ram_buffer(1234) := X"28AD000A";
		ram_buffer(1235) := X"11A00003";
		ram_buffer(1236) := X"00852021";
		ram_buffer(1237) := X"24040030";
		ram_buffer(1238) := X"00852021";
		ram_buffer(1239) := X"254A0001";
		ram_buffer(1240) := X"1120009F";
		ram_buffer(1241) := X"A1040000";
		ram_buffer(1242) := X"1000FFE6";
		ram_buffer(1243) := X"01604025";
		ram_buffer(1244) := X"8EB60000";
		ram_buffer(1245) := X"26B50004";
		ram_buffer(1246) := X"82C20000";
		ram_buffer(1247) := X"00000000";
		ram_buffer(1248) := X"104000ED";
		ram_buffer(1249) := X"26D40001";
		ram_buffer(1250) := X"12000018";
		ram_buffer(1251) := X"02802025";
		ram_buffer(1252) := X"10000004";
		ram_buffer(1253) := X"24840001";
		ram_buffer(1254) := X"10C00014";
		ram_buffer(1255) := X"00C08025";
		ram_buffer(1256) := X"24840001";
		ram_buffer(1257) := X"8085FFFF";
		ram_buffer(1258) := X"00000000";
		ram_buffer(1259) := X"14A0FFFA";
		ram_buffer(1260) := X"2606FFFF";
		ram_buffer(1261) := X"10C0000D";
		ram_buffer(1262) := X"2610FFFE";
		ram_buffer(1263) := X"060000D0";
		ram_buffer(1264) := X"00000000";
		ram_buffer(1265) := X"26100001";
		ram_buffer(1266) := X"00602025";
		ram_buffer(1267) := X"02003025";
		ram_buffer(1268) := X"0C000712";
		ram_buffer(1269) := X"24050020";
		ram_buffer(1270) := X"00401825";
		ram_buffer(1271) := X"82C20000";
		ram_buffer(1272) := X"00000000";
		ram_buffer(1273) := X"1040FEF7";
		ram_buffer(1274) := X"00701821";
		ram_buffer(1275) := X"24630001";
		ram_buffer(1276) := X"A062FFFF";
		ram_buffer(1277) := X"26940001";
		ram_buffer(1278) := X"8282FFFF";
		ram_buffer(1279) := X"00000000";
		ram_buffer(1280) := X"1040FEF0";
		ram_buffer(1281) := X"26940001";
		ram_buffer(1282) := X"24630001";
		ram_buffer(1283) := X"A062FFFF";
		ram_buffer(1284) := X"8282FFFF";
		ram_buffer(1285) := X"00000000";
		ram_buffer(1286) := X"1440FFF5";
		ram_buffer(1287) := X"24630001";
		ram_buffer(1288) := X"1000FEE8";
		ram_buffer(1289) := X"2463FFFF";
		ram_buffer(1290) := X"1482FEE6";
		ram_buffer(1291) := X"00000000";
		ram_buffer(1292) := X"8EA50000";
		ram_buffer(1293) := X"00000000";
		ram_buffer(1294) := X"2CA20010";
		ram_buffer(1295) := X"144000BA";
		ram_buffer(1296) := X"26B50004";
		ram_buffer(1297) := X"24020001";
		ram_buffer(1298) := X"00021100";
		ram_buffer(1299) := X"14400002";
		ram_buffer(1300) := X"00A2001B";
		ram_buffer(1301) := X"0007000D";
		ram_buffer(1302) := X"00003012";
		ram_buffer(1303) := X"2CC60010";
		ram_buffer(1304) := X"10C0FFF9";
		ram_buffer(1305) := X"00000000";
		ram_buffer(1306) := X"1040009D";
		ram_buffer(1307) := X"00000000";
		ram_buffer(1308) := X"24060058";
		ram_buffer(1309) := X"27A90010";
		ram_buffer(1310) := X"10860019";
		ram_buffer(1311) := X"00005025";
		ram_buffer(1312) := X"14400002";
		ram_buffer(1313) := X"00A2001B";
		ram_buffer(1314) := X"0007000D";
		ram_buffer(1315) := X"00002810";
		ram_buffer(1316) := X"00004012";
		ram_buffer(1317) := X"15400003";
		ram_buffer(1318) := X"00021102";
		ram_buffer(1319) := X"19000080";
		ram_buffer(1320) := X"00000000";
		ram_buffer(1321) := X"290B000A";
		ram_buffer(1322) := X"25240001";
		ram_buffer(1323) := X"11600002";
		ram_buffer(1324) := X"24060057";
		ram_buffer(1325) := X"24060030";
		ram_buffer(1326) := X"00C83021";
		ram_buffer(1327) := X"254A0001";
		ram_buffer(1328) := X"10400019";
		ram_buffer(1329) := X"A1260000";
		ram_buffer(1330) := X"1000FFED";
		ram_buffer(1331) := X"00804825";
		ram_buffer(1332) := X"10400076";
		ram_buffer(1333) := X"25060030";
		ram_buffer(1334) := X"01202025";
		ram_buffer(1335) := X"00804825";
		ram_buffer(1336) := X"14400002";
		ram_buffer(1337) := X"00A2001B";
		ram_buffer(1338) := X"0007000D";
		ram_buffer(1339) := X"00002810";
		ram_buffer(1340) := X"00004012";
		ram_buffer(1341) := X"15400003";
		ram_buffer(1342) := X"00021102";
		ram_buffer(1343) := X"1900FFF4";
		ram_buffer(1344) := X"00000000";
		ram_buffer(1345) := X"290B000A";
		ram_buffer(1346) := X"25240001";
		ram_buffer(1347) := X"11600002";
		ram_buffer(1348) := X"24060037";
		ram_buffer(1349) := X"24060030";
		ram_buffer(1350) := X"00C83021";
		ram_buffer(1351) := X"254A0001";
		ram_buffer(1352) := X"1440FFEE";
		ram_buffer(1353) := X"A1260000";
		ram_buffer(1354) := X"14E0002B";
		ram_buffer(1355) := X"A0800000";
		ram_buffer(1356) := X"24050020";
		ram_buffer(1357) := X"83B40010";
		ram_buffer(1358) := X"00000000";
		ram_buffer(1359) := X"1280006A";
		ram_buffer(1360) := X"00000000";
		ram_buffer(1361) := X"12000013";
		ram_buffer(1362) := X"27A20011";
		ram_buffer(1363) := X"10000004";
		ram_buffer(1364) := X"24420001";
		ram_buffer(1365) := X"10C0000F";
		ram_buffer(1366) := X"00C08025";
		ram_buffer(1367) := X"24420001";
		ram_buffer(1368) := X"8044FFFF";
		ram_buffer(1369) := X"00000000";
		ram_buffer(1370) := X"1480FFFA";
		ram_buffer(1371) := X"2606FFFF";
		ram_buffer(1372) := X"10C00008";
		ram_buffer(1373) := X"2610FFFE";
		ram_buffer(1374) := X"06000063";
		ram_buffer(1375) := X"00000000";
		ram_buffer(1376) := X"26100001";
		ram_buffer(1377) := X"00602025";
		ram_buffer(1378) := X"0C000712";
		ram_buffer(1379) := X"02003025";
		ram_buffer(1380) := X"00501821";
		ram_buffer(1381) := X"27A20011";
		ram_buffer(1382) := X"24630001";
		ram_buffer(1383) := X"24420001";
		ram_buffer(1384) := X"A074FFFF";
		ram_buffer(1385) := X"8054FFFF";
		ram_buffer(1386) := X"00000000";
		ram_buffer(1387) := X"1680FFFB";
		ram_buffer(1388) := X"24630001";
		ram_buffer(1389) := X"1000FE83";
		ram_buffer(1390) := X"2463FFFF";
		ram_buffer(1391) := X"A0720000";
		ram_buffer(1392) := X"1000FE80";
		ram_buffer(1393) := X"24630001";
		ram_buffer(1394) := X"1000FEC0";
		ram_buffer(1395) := X"01604025";
		ram_buffer(1396) := X"1000FEF8";
		ram_buffer(1397) := X"24050030";
		ram_buffer(1398) := X"1000FFD6";
		ram_buffer(1399) := X"24050030";
		ram_buffer(1400) := X"10E0002D";
		ram_buffer(1401) := X"A1600000";
		ram_buffer(1402) := X"24050030";
		ram_buffer(1403) := X"83B40010";
		ram_buffer(1404) := X"00000000";
		ram_buffer(1405) := X"1280003C";
		ram_buffer(1406) := X"00000000";
		ram_buffer(1407) := X"12000013";
		ram_buffer(1408) := X"27A20011";
		ram_buffer(1409) := X"10000004";
		ram_buffer(1410) := X"24420001";
		ram_buffer(1411) := X"10C0000F";
		ram_buffer(1412) := X"00C08025";
		ram_buffer(1413) := X"24420001";
		ram_buffer(1414) := X"8044FFFF";
		ram_buffer(1415) := X"00000000";
		ram_buffer(1416) := X"1480FFFA";
		ram_buffer(1417) := X"2606FFFF";
		ram_buffer(1418) := X"10C00008";
		ram_buffer(1419) := X"2610FFFE";
		ram_buffer(1420) := X"06000039";
		ram_buffer(1421) := X"00000000";
		ram_buffer(1422) := X"26100001";
		ram_buffer(1423) := X"00602025";
		ram_buffer(1424) := X"0C000712";
		ram_buffer(1425) := X"02003025";
		ram_buffer(1426) := X"00501821";
		ram_buffer(1427) := X"27A20011";
		ram_buffer(1428) := X"24630001";
		ram_buffer(1429) := X"24420001";
		ram_buffer(1430) := X"A074FFFF";
		ram_buffer(1431) := X"8054FFFF";
		ram_buffer(1432) := X"00000000";
		ram_buffer(1433) := X"1680FFFB";
		ram_buffer(1434) := X"24630001";
		ram_buffer(1435) := X"1000FE55";
		ram_buffer(1436) := X"2463FFFF";
		ram_buffer(1437) := X"11200004";
		ram_buffer(1438) := X"24A40030";
		ram_buffer(1439) := X"01005825";
		ram_buffer(1440) := X"1000FF20";
		ram_buffer(1441) := X"01604025";
		ram_buffer(1442) := X"250B0001";
		ram_buffer(1443) := X"A1040000";
		ram_buffer(1444) := X"14E0FFD5";
		ram_buffer(1445) := X"A1600000";
		ram_buffer(1446) := X"1000FFD4";
		ram_buffer(1447) := X"24050020";
		ram_buffer(1448) := X"14400008";
		ram_buffer(1449) := X"01202025";
		ram_buffer(1450) := X"25060030";
		ram_buffer(1451) := X"25240001";
		ram_buffer(1452) := X"A1260000";
		ram_buffer(1453) := X"10E0FF9E";
		ram_buffer(1454) := X"A0800000";
		ram_buffer(1455) := X"1000FF9D";
		ram_buffer(1456) := X"24050030";
		ram_buffer(1457) := X"1000FF6E";
		ram_buffer(1458) := X"00804825";
		ram_buffer(1459) := X"2402002D";
		ram_buffer(1460) := X"00052823";
		ram_buffer(1461) := X"A3A20010";
		ram_buffer(1462) := X"1000FEF8";
		ram_buffer(1463) := X"27A80011";
		ram_buffer(1464) := X"1000FF91";
		ram_buffer(1465) := X"27A40010";
		ram_buffer(1466) := X"1200FE36";
		ram_buffer(1467) := X"00602025";
		ram_buffer(1468) := X"0C000712";
		ram_buffer(1469) := X"02003025";
		ram_buffer(1470) := X"1000FE32";
		ram_buffer(1471) := X"00501821";
		ram_buffer(1472) := X"1000FF30";
		ram_buffer(1473) := X"00008025";
		ram_buffer(1474) := X"1000FF9D";
		ram_buffer(1475) := X"00008025";
		ram_buffer(1476) := X"1000FEBB";
		ram_buffer(1477) := X"00008025";
		ram_buffer(1478) := X"1000FFC7";
		ram_buffer(1479) := X"00008025";
		ram_buffer(1480) := X"1000FEF6";
		ram_buffer(1481) := X"24020001";
		ram_buffer(1482) := X"1000FF51";
		ram_buffer(1483) := X"24020001";
		ram_buffer(1484) := X"1000FE63";
		ram_buffer(1485) := X"24020001";
		ram_buffer(1486) := X"1200FE22";
		ram_buffer(1487) := X"2610FFFF";
		ram_buffer(1488) := X"1000FF1E";
		ram_buffer(1489) := X"00000000";
		ram_buffer(1490) := X"27BDFFE0";
		ram_buffer(1491) := X"AFBF001C";
		ram_buffer(1492) := X"AFB10018";
		ram_buffer(1493) := X"AFB00014";
		ram_buffer(1494) := X"3C111000";
		ram_buffer(1495) := X"8E222714";
		ram_buffer(1496) := X"00000000";
		ram_buffer(1497) := X"8C420004";
		ram_buffer(1498) := X"00000000";
		ram_buffer(1499) := X"2C430008";
		ram_buffer(1500) := X"1060000F";
		ram_buffer(1501) := X"3C101000";
		ram_buffer(1502) := X"26102718";
		ram_buffer(1503) := X"000210C0";
		ram_buffer(1504) := X"02021021";
		ram_buffer(1505) := X"8C430000";
		ram_buffer(1506) := X"8C440004";
		ram_buffer(1507) := X"0060F809";
		ram_buffer(1508) := X"00000000";
		ram_buffer(1509) := X"8E222714";
		ram_buffer(1510) := X"00000000";
		ram_buffer(1511) := X"8C420004";
		ram_buffer(1512) := X"00000000";
		ram_buffer(1513) := X"2C430008";
		ram_buffer(1514) := X"1460FFF4";
		ram_buffer(1515) := X"00000000";
		ram_buffer(1516) := X"8FBF001C";
		ram_buffer(1517) := X"8FB10018";
		ram_buffer(1518) := X"8FB00014";
		ram_buffer(1519) := X"03E00008";
		ram_buffer(1520) := X"27BD0020";
		ram_buffer(1521) := X"8F828018";
		ram_buffer(1522) := X"00000000";
		ram_buffer(1523) := X"8C430004";
		ram_buffer(1524) := X"8F828010";
		ram_buffer(1525) := X"8F84800C";
		ram_buffer(1526) := X"24420001";
		ram_buffer(1527) := X"304201FF";
		ram_buffer(1528) := X"10440008";
		ram_buffer(1529) := X"00000000";
		ram_buffer(1530) := X"8F848010";
		ram_buffer(1531) := X"3C051000";
		ram_buffer(1532) := X"24A52508";
		ram_buffer(1533) := X"306300FF";
		ram_buffer(1534) := X"00852021";
		ram_buffer(1535) := X"A0830000";
		ram_buffer(1536) := X"AF828010";
		ram_buffer(1537) := X"03E00008";
		ram_buffer(1538) := X"00000000";
		ram_buffer(1539) := X"3C02F000";
		ram_buffer(1540) := X"8C430004";
		ram_buffer(1541) := X"3C021000";
		ram_buffer(1542) := X"00032080";
		ram_buffer(1543) := X"24422708";
		ram_buffer(1544) := X"00441021";
		ram_buffer(1545) := X"3C031000";
		ram_buffer(1546) := X"24632758";
		ram_buffer(1547) := X"00641821";
		ram_buffer(1548) := X"8C630000";
		ram_buffer(1549) := X"24040007";
		ram_buffer(1550) := X"AC640000";
		ram_buffer(1551) := X"8C430000";
		ram_buffer(1552) := X"00000000";
		ram_buffer(1553) := X"24630001";
		ram_buffer(1554) := X"03E00008";
		ram_buffer(1555) := X"AC430000";
		ram_buffer(1556) := X"8F838018";
		ram_buffer(1557) := X"00000000";
		ram_buffer(1558) := X"8C620000";
		ram_buffer(1559) := X"00000000";
		ram_buffer(1560) := X"30420002";
		ram_buffer(1561) := X"1040FFFC";
		ram_buffer(1562) := X"00000000";
		ram_buffer(1563) := X"AC650008";
		ram_buffer(1564) := X"03E00008";
		ram_buffer(1565) := X"00000000";
		ram_buffer(1566) := X"3C022000";
		ram_buffer(1567) := X"AF82801C";
		ram_buffer(1568) := X"3C051000";
		ram_buffer(1569) := X"3C022004";
		ram_buffer(1570) := X"27BDFFE8";
		ram_buffer(1571) := X"AF828018";
		ram_buffer(1572) := X"24A51850";
		ram_buffer(1573) := X"3C022003";
		ram_buffer(1574) := X"AF828014";
		ram_buffer(1575) := X"AFBF0014";
		ram_buffer(1576) := X"0C0003CD";
		ram_buffer(1577) := X"00002025";
		ram_buffer(1578) := X"3C041000";
		ram_buffer(1579) := X"3C032001";
		ram_buffer(1580) := X"AC832714";
		ram_buffer(1581) := X"3C031000";
		ram_buffer(1582) := X"24822714";
		ram_buffer(1583) := X"246317C4";
		ram_buffer(1584) := X"AC400004";
		ram_buffer(1585) := X"AC40000C";
		ram_buffer(1586) := X"AC40001C";
		ram_buffer(1587) := X"AC400024";
		ram_buffer(1588) := X"AC40002C";
		ram_buffer(1589) := X"AC400034";
		ram_buffer(1590) := X"AC40003C";
		ram_buffer(1591) := X"AC430014";
		ram_buffer(1592) := X"AC400018";
		ram_buffer(1593) := X"3C06F000";
		ram_buffer(1594) := X"8CC30004";
		ram_buffer(1595) := X"3C051000";
		ram_buffer(1596) := X"00031100";
		ram_buffer(1597) := X"00431021";
		ram_buffer(1598) := X"00021080";
		ram_buffer(1599) := X"3C031000";
		ram_buffer(1600) := X"24631D98";
		ram_buffer(1601) := X"24420004";
		ram_buffer(1602) := X"00621021";
		ram_buffer(1603) := X"24A51748";
		ram_buffer(1604) := X"AC450038";
		ram_buffer(1605) := X"AC40003C";
		ram_buffer(1606) := X"8CC50004";
		ram_buffer(1607) := X"00000000";
		ram_buffer(1608) := X"00051100";
		ram_buffer(1609) := X"00451021";
		ram_buffer(1610) := X"00021080";
		ram_buffer(1611) := X"00431021";
		ram_buffer(1612) := X"8C420000";
		ram_buffer(1613) := X"24030082";
		ram_buffer(1614) := X"AC430000";
		ram_buffer(1615) := X"8C822714";
		ram_buffer(1616) := X"8FBF0014";
		ram_buffer(1617) := X"24030005";
		ram_buffer(1618) := X"AC430000";
		ram_buffer(1619) := X"08000049";
		ram_buffer(1620) := X"27BD0018";
		ram_buffer(1621) := X"3C06F000";
		ram_buffer(1622) := X"8CC70004";
		ram_buffer(1623) := X"3C031000";
		ram_buffer(1624) := X"00071080";
		ram_buffer(1625) := X"24632758";
		ram_buffer(1626) := X"00621821";
		ram_buffer(1627) := X"3C02F003";
		ram_buffer(1628) := X"AC620000";
		ram_buffer(1629) := X"8C620000";
		ram_buffer(1630) := X"3404C350";
		ram_buffer(1631) := X"AC440004";
		ram_buffer(1632) := X"8CC40004";
		ram_buffer(1633) := X"3C051000";
		ram_buffer(1634) := X"00041100";
		ram_buffer(1635) := X"00441021";
		ram_buffer(1636) := X"00021080";
		ram_buffer(1637) := X"3C041000";
		ram_buffer(1638) := X"24420004";
		ram_buffer(1639) := X"24841D98";
		ram_buffer(1640) := X"00821021";
		ram_buffer(1641) := X"24A5180C";
		ram_buffer(1642) := X"AC450008";
		ram_buffer(1643) := X"10E0000A";
		ram_buffer(1644) := X"AC40000C";
		ram_buffer(1645) := X"8CC50004";
		ram_buffer(1646) := X"00000000";
		ram_buffer(1647) := X"00051100";
		ram_buffer(1648) := X"00451021";
		ram_buffer(1649) := X"00021080";
		ram_buffer(1650) := X"00441021";
		ram_buffer(1651) := X"8C420000";
		ram_buffer(1652) := X"24040002";
		ram_buffer(1653) := X"AC440000";
		ram_buffer(1654) := X"8C620000";
		ram_buffer(1655) := X"24030003";
		ram_buffer(1656) := X"AC430000";
		ram_buffer(1657) := X"08000046";
		ram_buffer(1658) := X"24040001";
		ram_buffer(1659) := X"8F838018";
		ram_buffer(1660) := X"00000000";
		ram_buffer(1661) := X"8C620000";
		ram_buffer(1662) := X"00000000";
		ram_buffer(1663) := X"30420002";
		ram_buffer(1664) := X"1040FFFC";
		ram_buffer(1665) := X"00000000";
		ram_buffer(1666) := X"AC640008";
		ram_buffer(1667) := X"03E00008";
		ram_buffer(1668) := X"00000000";
		ram_buffer(1669) := X"10000003";
		ram_buffer(1670) := X"00000000";
		ram_buffer(1671) := X"40836000";
		ram_buffer(1672) := X"00000000";
		ram_buffer(1673) := X"40036000";
		ram_buffer(1674) := X"40806000";
		ram_buffer(1675) := X"8F848010";
		ram_buffer(1676) := X"8F82800C";
		ram_buffer(1677) := X"00000000";
		ram_buffer(1678) := X"1082FFF8";
		ram_buffer(1679) := X"00000000";
		ram_buffer(1680) := X"8F82800C";
		ram_buffer(1681) := X"3C041000";
		ram_buffer(1682) := X"24842508";
		ram_buffer(1683) := X"00441021";
		ram_buffer(1684) := X"90420000";
		ram_buffer(1685) := X"8F84800C";
		ram_buffer(1686) := X"304200FF";
		ram_buffer(1687) := X"24840001";
		ram_buffer(1688) := X"308401FF";
		ram_buffer(1689) := X"AF84800C";
		ram_buffer(1690) := X"40836000";
		ram_buffer(1691) := X"03E00008";
		ram_buffer(1692) := X"00000000";
		ram_buffer(1693) := X"24050004";
		ram_buffer(1694) := X"8F838018";
		ram_buffer(1695) := X"308600FF";
		ram_buffer(1696) := X"8C620000";
		ram_buffer(1697) := X"00000000";
		ram_buffer(1698) := X"30420002";
		ram_buffer(1699) := X"1040FFFC";
		ram_buffer(1700) := X"00000000";
		ram_buffer(1701) := X"24A5FFFF";
		ram_buffer(1702) := X"AC660008";
		ram_buffer(1703) := X"14A0FFF6";
		ram_buffer(1704) := X"00042202";
		ram_buffer(1705) := X"03E00008";
		ram_buffer(1706) := X"00000000";
		ram_buffer(1707) := X"3C071000";
		ram_buffer(1708) := X"00003025";
		ram_buffer(1709) := X"00001025";
		ram_buffer(1710) := X"24E72508";
		ram_buffer(1711) := X"24080020";
		ram_buffer(1712) := X"40036000";
		ram_buffer(1713) := X"40806000";
		ram_buffer(1714) := X"8F858010";
		ram_buffer(1715) := X"8F84800C";
		ram_buffer(1716) := X"00000000";
		ram_buffer(1717) := X"14A4000A";
		ram_buffer(1718) := X"00000000";
		ram_buffer(1719) := X"40836000";
		ram_buffer(1720) := X"00000000";
		ram_buffer(1721) := X"40036000";
		ram_buffer(1722) := X"40806000";
		ram_buffer(1723) := X"8F858010";
		ram_buffer(1724) := X"8F84800C";
		ram_buffer(1725) := X"00000000";
		ram_buffer(1726) := X"10A4FFF8";
		ram_buffer(1727) := X"00000000";
		ram_buffer(1728) := X"8F84800C";
		ram_buffer(1729) := X"00000000";
		ram_buffer(1730) := X"00E42021";
		ram_buffer(1731) := X"90840000";
		ram_buffer(1732) := X"8F85800C";
		ram_buffer(1733) := X"308400FF";
		ram_buffer(1734) := X"24A50001";
		ram_buffer(1735) := X"30A501FF";
		ram_buffer(1736) := X"AF85800C";
		ram_buffer(1737) := X"40836000";
		ram_buffer(1738) := X"00C41804";
		ram_buffer(1739) := X"24C60008";
		ram_buffer(1740) := X"14C8FFE3";
		ram_buffer(1741) := X"00431025";
		ram_buffer(1742) := X"03E00008";
		ram_buffer(1743) := X"00000000";
		ram_buffer(1744) := X"8F828014";
		ram_buffer(1745) := X"00000000";
		ram_buffer(1746) := X"03E00008";
		ram_buffer(1747) := X"AC440008";
		ram_buffer(1748) := X"8F828014";
		ram_buffer(1749) := X"00000000";
		ram_buffer(1750) := X"8C420008";
		ram_buffer(1751) := X"03E00008";
		ram_buffer(1752) := X"00000000";
		ram_buffer(1753) := X"8F828014";
		ram_buffer(1754) := X"00000000";
		ram_buffer(1755) := X"8C420004";
		ram_buffer(1756) := X"03E00008";
		ram_buffer(1757) := X"00000000";
		ram_buffer(1758) := X"3C03F000";
		ram_buffer(1759) := X"8C620004";
		ram_buffer(1760) := X"00000000";
		ram_buffer(1761) := X"24420001";
		ram_buffer(1762) := X"8F84801C";
		ram_buffer(1763) := X"00000000";
		ram_buffer(1764) := X"AC820000";
		ram_buffer(1765) := X"8C620004";
		ram_buffer(1766) := X"8F84801C";
		ram_buffer(1767) := X"24420001";
		ram_buffer(1768) := X"8C840000";
		ram_buffer(1769) := X"00000000";
		ram_buffer(1770) := X"1444FFF4";
		ram_buffer(1771) := X"00000000";
		ram_buffer(1772) := X"080001AD";
		ram_buffer(1773) := X"00000000";
		ram_buffer(1774) := X"27BDFFE8";
		ram_buffer(1775) := X"AFBF0014";
		ram_buffer(1776) := X"0C0001AD";
		ram_buffer(1777) := X"00000000";
		ram_buffer(1778) := X"3C02F000";
		ram_buffer(1779) := X"8C420004";
		ram_buffer(1780) := X"00000000";
		ram_buffer(1781) := X"24420001";
		ram_buffer(1782) := X"8FBF0014";
		ram_buffer(1783) := X"8F83801C";
		ram_buffer(1784) := X"00000000";
		ram_buffer(1785) := X"AC620000";
		ram_buffer(1786) := X"03E00008";
		ram_buffer(1787) := X"27BD0018";
		ram_buffer(1788) := X"3C031000";
		ram_buffer(1789) := X"24632708";
		ram_buffer(1790) := X"3C05F000";
		ram_buffer(1791) := X"8CA20004";
		ram_buffer(1792) := X"00000000";
		ram_buffer(1793) := X"00021080";
		ram_buffer(1794) := X"00621021";
		ram_buffer(1795) := X"8C420000";
		ram_buffer(1796) := X"00000000";
		ram_buffer(1797) := X"1482FFF9";
		ram_buffer(1798) := X"00000000";
		ram_buffer(1799) := X"03E00008";
		ram_buffer(1800) := X"00000000";
		ram_buffer(1801) := X"3C02F000";
		ram_buffer(1802) := X"8C420004";
		ram_buffer(1803) := X"3C031000";
		ram_buffer(1804) := X"24632708";
		ram_buffer(1805) := X"00021080";
		ram_buffer(1806) := X"00431021";
		ram_buffer(1807) := X"8C420000";
		ram_buffer(1808) := X"03E00008";
		ram_buffer(1809) := X"00000000";
		ram_buffer(1810) := X"28CA0008";
		ram_buffer(1811) := X"1540003E";
		ram_buffer(1812) := X"00801025";
		ram_buffer(1813) := X"10A00007";
		ram_buffer(1814) := X"00043823";
		ram_buffer(1815) := X"00000000";
		ram_buffer(1816) := X"30A500FF";
		ram_buffer(1817) := X"00055200";
		ram_buffer(1818) := X"00AA2825";
		ram_buffer(1819) := X"00055400";
		ram_buffer(1820) := X"00AA2825";
		ram_buffer(1821) := X"30EA0003";
		ram_buffer(1822) := X"11400003";
		ram_buffer(1823) := X"00CA3023";
		ram_buffer(1824) := X"A8850000";
		ram_buffer(1825) := X"008A2021";
		ram_buffer(1826) := X"30EA0004";
		ram_buffer(1827) := X"11400003";
		ram_buffer(1828) := X"00CA3023";
		ram_buffer(1829) := X"AC850000";
		ram_buffer(1830) := X"008A2021";
		ram_buffer(1831) := X"30D8003F";
		ram_buffer(1832) := X"10D80016";
		ram_buffer(1833) := X"00D83823";
		ram_buffer(1834) := X"00873821";
		ram_buffer(1835) := X"AC850000";
		ram_buffer(1836) := X"AC850004";
		ram_buffer(1837) := X"AC850008";
		ram_buffer(1838) := X"AC85000C";
		ram_buffer(1839) := X"AC850010";
		ram_buffer(1840) := X"AC850014";
		ram_buffer(1841) := X"AC850018";
		ram_buffer(1842) := X"AC85001C";
		ram_buffer(1843) := X"AC850020";
		ram_buffer(1844) := X"AC850024";
		ram_buffer(1845) := X"AC850028";
		ram_buffer(1846) := X"AC85002C";
		ram_buffer(1847) := X"AC850030";
		ram_buffer(1848) := X"AC850034";
		ram_buffer(1849) := X"AC850038";
		ram_buffer(1850) := X"AC85003C";
		ram_buffer(1851) := X"24840040";
		ram_buffer(1852) := X"1487FFEE";
		ram_buffer(1853) := X"00000000";
		ram_buffer(1854) := X"03003025";
		ram_buffer(1855) := X"30D8001F";
		ram_buffer(1856) := X"10D8000A";
		ram_buffer(1857) := X"00000000";
		ram_buffer(1858) := X"AC850000";
		ram_buffer(1859) := X"AC850004";
		ram_buffer(1860) := X"AC850008";
		ram_buffer(1861) := X"AC85000C";
		ram_buffer(1862) := X"AC850010";
		ram_buffer(1863) := X"AC850014";
		ram_buffer(1864) := X"AC850018";
		ram_buffer(1865) := X"AC85001C";
		ram_buffer(1866) := X"24840020";
		ram_buffer(1867) := X"33060003";
		ram_buffer(1868) := X"10D80005";
		ram_buffer(1869) := X"03063823";
		ram_buffer(1870) := X"00873821";
		ram_buffer(1871) := X"24840004";
		ram_buffer(1872) := X"1487FFFE";
		ram_buffer(1873) := X"AC85FFFC";
		ram_buffer(1874) := X"18C00004";
		ram_buffer(1875) := X"00863821";
		ram_buffer(1876) := X"24840001";
		ram_buffer(1877) := X"1487FFFE";
		ram_buffer(1878) := X"A085FFFF";
		ram_buffer(1879) := X"03E00008";
		ram_buffer(1880) := X"00000000";
		ram_buffer(1881) := X"00000000";
		ram_buffer(1882) := X"00000100";
		ram_buffer(1883) := X"01010001";
		ram_buffer(1884) := X"00000000";
		ram_buffer(1885) := X"00000000";
		ram_buffer(1886) := X"00000000";
		ram_buffer(1887) := X"00000000";
		ram_buffer(1888) := X"FFFFFFFF";
		ram_buffer(1889) := X"FFFFFFFF";
		ram_buffer(1890) := X"FFFFFFFF";
		ram_buffer(1891) := X"FFFFFFFF";
		ram_buffer(1892) := X"FFFFFFFF";
		ram_buffer(1893) := X"FFFFFFFF";
		ram_buffer(1894) := X"FFFFFFFF";
		ram_buffer(1895) := X"00000000";
		ram_buffer(1896) := X"00000000";
		ram_buffer(1897) := X"00000000";
		ram_buffer(1898) := X"00000000";
		ram_buffer(1899) := X"00000000";
		ram_buffer(1900) := X"00000000";
		ram_buffer(1901) := X"00000000";
		ram_buffer(1902) := X"00000000";
		ram_buffer(1903) := X"00000000";
		ram_buffer(1904) := X"00000000";
		ram_buffer(1905) := X"00000000";
		ram_buffer(1906) := X"00000000";
		ram_buffer(1907) := X"00000000";
		ram_buffer(1908) := X"00000000";
		ram_buffer(1909) := X"00000000";
		ram_buffer(1910) := X"00000000";
		ram_buffer(1911) := X"FFFFFFFF";
		ram_buffer(1912) := X"00000000";
		ram_buffer(1913) := X"00000000";
		ram_buffer(1914) := X"00000000";
		ram_buffer(1915) := X"00000000";
		ram_buffer(1916) := X"00000000";
		ram_buffer(1917) := X"00000000";
		ram_buffer(1918) := X"00000000";
		ram_buffer(1919) := X"00000000";
		ram_buffer(1920) := X"00000000";
		ram_buffer(1921) := X"00000000";
		ram_buffer(1922) := X"00000000";
		ram_buffer(1923) := X"00000000";
		ram_buffer(1924) := X"00000000";
		ram_buffer(1925) := X"00000000";
		ram_buffer(1926) := X"00000000";
		ram_buffer(1927) := X"00000000";
		ram_buffer(1928) := X"FFFFFFFF";
		ram_buffer(1929) := X"00000000";
		ram_buffer(1930) := X"00000000";
		ram_buffer(1931) := X"00000000";
		ram_buffer(1932) := X"00000000";
		ram_buffer(1933) := X"00000000";
		ram_buffer(1934) := X"00000000";
		ram_buffer(1935) := X"00000000";
		ram_buffer(1936) := X"00000000";
		ram_buffer(1937) := X"00000000";
		ram_buffer(1938) := X"00000000";
		ram_buffer(1939) := X"00000000";
		ram_buffer(1940) := X"00000000";
		ram_buffer(1941) := X"00000000";
		ram_buffer(1942) := X"00000000";
		ram_buffer(1943) := X"00000000";
		ram_buffer(1944) := X"00000000";
		return ram_buffer;
	end;
end;
