library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

package koc_lock_pack is
    constant axi_resp_okay : std_logic_vector := "00";
end package;