library ieee;
use ieee.std_logic_1164.all;

package main_pack is

	constant cpu_width : integer := 32;
	constant ram_size : integer := 1003;
	subtype word_type is std_logic_vector(cpu_width-1 downto 0);
	type ram_type is array(0 to ram_size-1) of word_type;
	function load_hex return ram_type;

end package;

package body main_pack is

	function load_hex return ram_type is
		variable ram_buffer : ram_type := (others=>(others=>'0'));
	begin
		ram_buffer(0) := X"3C1C1001";
		ram_buffer(1) := X"279C8FA0";
		ram_buffer(2) := X"3C1D1000";
		ram_buffer(3) := X"27BD0FE8";
		ram_buffer(4) := X"0C0000E0";
		ram_buffer(5) := X"00000000";
		ram_buffer(6) := X"00000000";
		ram_buffer(7) := X"00000000";
		ram_buffer(8) := X"00000000";
		ram_buffer(9) := X"00000000";
		ram_buffer(10) := X"00000000";
		ram_buffer(11) := X"00000000";
		ram_buffer(12) := X"00000000";
		ram_buffer(13) := X"00000000";
		ram_buffer(14) := X"00000000";
		ram_buffer(15) := X"23BDFF98";
		ram_buffer(16) := X"AFA10010";
		ram_buffer(17) := X"AFA20014";
		ram_buffer(18) := X"AFA30018";
		ram_buffer(19) := X"AFA4001C";
		ram_buffer(20) := X"AFA50020";
		ram_buffer(21) := X"AFA60024";
		ram_buffer(22) := X"AFA70028";
		ram_buffer(23) := X"AFA8002C";
		ram_buffer(24) := X"AFA90030";
		ram_buffer(25) := X"AFAA0034";
		ram_buffer(26) := X"AFAB0038";
		ram_buffer(27) := X"AFAC003C";
		ram_buffer(28) := X"AFAD0040";
		ram_buffer(29) := X"AFAE0044";
		ram_buffer(30) := X"AFAF0048";
		ram_buffer(31) := X"AFB8004C";
		ram_buffer(32) := X"AFB90050";
		ram_buffer(33) := X"AFBF0054";
		ram_buffer(34) := X"401A7000";
		ram_buffer(35) := X"235AFFFC";
		ram_buffer(36) := X"AFBA0058";
		ram_buffer(37) := X"0000D810";
		ram_buffer(38) := X"AFBB005C";
		ram_buffer(39) := X"0000D812";
		ram_buffer(40) := X"AFBB0060";
		ram_buffer(41) := X"0C0000B8";
		ram_buffer(42) := X"23A50000";
		ram_buffer(43) := X"8FA10010";
		ram_buffer(44) := X"8FA20014";
		ram_buffer(45) := X"8FA30018";
		ram_buffer(46) := X"8FA4001C";
		ram_buffer(47) := X"8FA50020";
		ram_buffer(48) := X"8FA60024";
		ram_buffer(49) := X"8FA70028";
		ram_buffer(50) := X"8FA8002C";
		ram_buffer(51) := X"8FA90030";
		ram_buffer(52) := X"8FAA0034";
		ram_buffer(53) := X"8FAB0038";
		ram_buffer(54) := X"8FAC003C";
		ram_buffer(55) := X"8FAD0040";
		ram_buffer(56) := X"8FAE0044";
		ram_buffer(57) := X"8FAF0048";
		ram_buffer(58) := X"8FB8004C";
		ram_buffer(59) := X"8FB90050";
		ram_buffer(60) := X"8FBF0054";
		ram_buffer(61) := X"8FBA0058";
		ram_buffer(62) := X"8FBB005C";
		ram_buffer(63) := X"03600011";
		ram_buffer(64) := X"8FBB0060";
		ram_buffer(65) := X"03600013";
		ram_buffer(66) := X"23BD0068";
		ram_buffer(67) := X"341B0001";
		ram_buffer(68) := X"03400008";
		ram_buffer(69) := X"409B6000";
		ram_buffer(70) := X"40026000";
		ram_buffer(71) := X"03E00008";
		ram_buffer(72) := X"40846000";
		ram_buffer(73) := X"3C051000";
		ram_buffer(74) := X"24A50150";
		ram_buffer(75) := X"8CA60000";
		ram_buffer(76) := X"AC06003C";
		ram_buffer(77) := X"8CA60004";
		ram_buffer(78) := X"AC060040";
		ram_buffer(79) := X"8CA60008";
		ram_buffer(80) := X"AC060044";
		ram_buffer(81) := X"8CA6000C";
		ram_buffer(82) := X"03E00008";
		ram_buffer(83) := X"AC060048";
		ram_buffer(84) := X"3C1A1000";
		ram_buffer(85) := X"375A003C";
		ram_buffer(86) := X"03400008";
		ram_buffer(87) := X"00000000";
		ram_buffer(88) := X"00850019";
		ram_buffer(89) := X"00001012";
		ram_buffer(90) := X"00002010";
		ram_buffer(91) := X"03E00008";
		ram_buffer(92) := X"ACC40000";
		ram_buffer(93) := X"0000000C";
		ram_buffer(94) := X"03E00008";
		ram_buffer(95) := X"00000000";
		ram_buffer(96) := X"AC900000";
		ram_buffer(97) := X"AC910004";
		ram_buffer(98) := X"AC920008";
		ram_buffer(99) := X"AC93000C";
		ram_buffer(100) := X"AC940010";
		ram_buffer(101) := X"AC950014";
		ram_buffer(102) := X"AC960018";
		ram_buffer(103) := X"AC97001C";
		ram_buffer(104) := X"AC9E0020";
		ram_buffer(105) := X"AC9C0024";
		ram_buffer(106) := X"AC9D0028";
		ram_buffer(107) := X"AC9F002C";
		ram_buffer(108) := X"03E00008";
		ram_buffer(109) := X"34020000";
		ram_buffer(110) := X"8C900000";
		ram_buffer(111) := X"8C910004";
		ram_buffer(112) := X"8C920008";
		ram_buffer(113) := X"8C93000C";
		ram_buffer(114) := X"8C940010";
		ram_buffer(115) := X"8C950014";
		ram_buffer(116) := X"8C960018";
		ram_buffer(117) := X"8C97001C";
		ram_buffer(118) := X"8C9E0020";
		ram_buffer(119) := X"8C9C0024";
		ram_buffer(120) := X"8C9D0028";
		ram_buffer(121) := X"8C9F002C";
		ram_buffer(122) := X"03E00008";
		ram_buffer(123) := X"34A20000";
		ram_buffer(124) := X"27BDFFE0";
		ram_buffer(125) := X"AFBF001C";
		ram_buffer(126) := X"AFB10018";
		ram_buffer(127) := X"0C0002B2";
		ram_buffer(128) := X"AFB00014";
		ram_buffer(129) := X"0C000391";
		ram_buffer(130) := X"24040001";
		ram_buffer(131) := X"3C101000";
		ram_buffer(132) := X"3C111000";
		ram_buffer(133) := X"3C051000";
		ram_buffer(134) := X"26100EC8";
		ram_buffer(135) := X"26310254";
		ram_buffer(136) := X"24060004";
		ram_buffer(137) := X"24A50ECC";
		ram_buffer(138) := X"24040004";
		ram_buffer(139) := X"0C000141";
		ram_buffer(140) := X"AE110004";
		ram_buffer(141) := X"3C051000";
		ram_buffer(142) := X"24060004";
		ram_buffer(143) := X"24A50ED0";
		ram_buffer(144) := X"24040004";
		ram_buffer(145) := X"0C000141";
		ram_buffer(146) := X"AE110008";
		ram_buffer(147) := X"0C000095";
		ram_buffer(148) := X"00000000";
		ram_buffer(149) := X"27BDFFE8";
		ram_buffer(150) := X"AFBF0014";
		ram_buffer(151) := X"0C000307";
		ram_buffer(152) := X"00000000";
		ram_buffer(153) := X"0C000395";
		ram_buffer(154) := X"00000000";
		ram_buffer(155) := X"2785800C";
		ram_buffer(156) := X"24060004";
		ram_buffer(157) := X"0C000141";
		ram_buffer(158) := X"00002025";
		ram_buffer(159) := X"8F84800C";
		ram_buffer(160) := X"0C000391";
		ram_buffer(161) := X"00000000";
		ram_buffer(162) := X"8F82800C";
		ram_buffer(163) := X"24060004";
		ram_buffer(164) := X"24420001";
		ram_buffer(165) := X"2785800C";
		ram_buffer(166) := X"24040004";
		ram_buffer(167) := X"AF82800C";
		ram_buffer(168) := X"0C000141";
		ram_buffer(169) := X"00000000";
		ram_buffer(170) := X"0C0003A4";
		ram_buffer(171) := X"00000000";
		ram_buffer(172) := X"1000FFEC";
		ram_buffer(173) := X"00000000";
		ram_buffer(174) := X"3C02F000";
		ram_buffer(175) := X"8C420004";
		ram_buffer(176) := X"3C031000";
		ram_buffer(177) := X"24630ED4";
		ram_buffer(178) := X"00021080";
		ram_buffer(179) := X"00431021";
		ram_buffer(180) := X"8C420000";
		ram_buffer(181) := X"24030002";
		ram_buffer(182) := X"03E00008";
		ram_buffer(183) := X"AC430000";
		ram_buffer(184) := X"27BDFFE0";
		ram_buffer(185) := X"AFBF001C";
		ram_buffer(186) := X"AFB20018";
		ram_buffer(187) := X"AFB10014";
		ram_buffer(188) := X"AFB00010";
		ram_buffer(189) := X"3C02F000";
		ram_buffer(190) := X"8C430004";
		ram_buffer(191) := X"00000000";
		ram_buffer(192) := X"00031100";
		ram_buffer(193) := X"00431021";
		ram_buffer(194) := X"00021080";
		ram_buffer(195) := X"24520004";
		ram_buffer(196) := X"3C111000";
		ram_buffer(197) := X"26310EE0";
		ram_buffer(198) := X"02221021";
		ram_buffer(199) := X"8C430000";
		ram_buffer(200) := X"00408025";
		ram_buffer(201) := X"8C630004";
		ram_buffer(202) := X"00000000";
		ram_buffer(203) := X"2C620008";
		ram_buffer(204) := X"14400007";
		ram_buffer(205) := X"00000000";
		ram_buffer(206) := X"8FBF001C";
		ram_buffer(207) := X"8FB20018";
		ram_buffer(208) := X"8FB10014";
		ram_buffer(209) := X"8FB00010";
		ram_buffer(210) := X"03E00008";
		ram_buffer(211) := X"27BD0020";
		ram_buffer(212) := X"000318C0";
		ram_buffer(213) := X"00721821";
		ram_buffer(214) := X"02231821";
		ram_buffer(215) := X"8C620000";
		ram_buffer(216) := X"8C640004";
		ram_buffer(217) := X"0040F809";
		ram_buffer(218) := X"00000000";
		ram_buffer(219) := X"8E020000";
		ram_buffer(220) := X"00000000";
		ram_buffer(221) := X"8C430004";
		ram_buffer(222) := X"1000FFED";
		ram_buffer(223) := X"2C620008";
		ram_buffer(224) := X"27BDFFD0";
		ram_buffer(225) := X"AFBF002C";
		ram_buffer(226) := X"AFB50028";
		ram_buffer(227) := X"AFB40024";
		ram_buffer(228) := X"AFB30020";
		ram_buffer(229) := X"AFB2001C";
		ram_buffer(230) := X"AFB10018";
		ram_buffer(231) := X"AFB00014";
		ram_buffer(232) := X"3C04F000";
		ram_buffer(233) := X"8C820004";
		ram_buffer(234) := X"00000000";
		ram_buffer(235) := X"00021240";
		ram_buffer(236) := X"244301E8";
		ram_buffer(237) := X"3C021000";
		ram_buffer(238) := X"24421000";
		ram_buffer(239) := X"00431021";
		ram_buffer(240) := X"0040E825";
		ram_buffer(241) := X"8C920004";
		ram_buffer(242) := X"8C950004";
		ram_buffer(243) := X"3C111000";
		ram_buffer(244) := X"00159900";
		ram_buffer(245) := X"02758021";
		ram_buffer(246) := X"00108080";
		ram_buffer(247) := X"26310EE0";
		ram_buffer(248) := X"0230A021";
		ram_buffer(249) := X"8C850004";
		ram_buffer(250) := X"3C021000";
		ram_buffer(251) := X"24420ED4";
		ram_buffer(252) := X"00052880";
		ram_buffer(253) := X"00A22821";
		ram_buffer(254) := X"3C02F002";
		ram_buffer(255) := X"ACA20000";
		ram_buffer(256) := X"24040004";
		ram_buffer(257) := X"0C000141";
		ram_buffer(258) := X"24060004";
		ram_buffer(259) := X"3C02F001";
		ram_buffer(260) := X"AE820000";
		ram_buffer(261) := X"26020004";
		ram_buffer(262) := X"02221021";
		ram_buffer(263) := X"26840044";
		ram_buffer(264) := X"00401825";
		ram_buffer(265) := X"14830020";
		ram_buffer(266) := X"24630008";
		ram_buffer(267) := X"3C031000";
		ram_buffer(268) := X"246302B8";
		ram_buffer(269) := X"AC430000";
		ram_buffer(270) := X"AC400004";
		ram_buffer(271) := X"02759821";
		ram_buffer(272) := X"00139880";
		ram_buffer(273) := X"02338821";
		ram_buffer(274) := X"8E220000";
		ram_buffer(275) := X"24030001";
		ram_buffer(276) := X"AC430000";
		ram_buffer(277) := X"24060004";
		ram_buffer(278) := X"02802825";
		ram_buffer(279) := X"0C000141";
		ram_buffer(280) := X"24040004";
		ram_buffer(281) := X"16400014";
		ram_buffer(282) := X"3C101000";
		ram_buffer(283) := X"2786800C";
		ram_buffer(284) := X"278288A4";
		ram_buffer(285) := X"14C2000E";
		ram_buffer(286) := X"24C60004";
		ram_buffer(287) := X"24C6FFFC";
		ram_buffer(288) := X"2782800C";
		ram_buffer(289) := X"24C60004";
		ram_buffer(290) := X"00C23023";
		ram_buffer(291) := X"00402825";
		ram_buffer(292) := X"0C000141";
		ram_buffer(293) := X"24040004";
		ram_buffer(294) := X"0C00007C";
		ram_buffer(295) := X"00000000";
		ram_buffer(296) := X"1000FFFF";
		ram_buffer(297) := X"00000000";
		ram_buffer(298) := X"1000FFDE";
		ram_buffer(299) := X"AC60FFF8";
		ram_buffer(300) := X"1000FFF0";
		ram_buffer(301) := X"ACC0FFFC";
		ram_buffer(302) := X"26100EC8";
		ram_buffer(303) := X"00129080";
		ram_buffer(304) := X"3C13F000";
		ram_buffer(305) := X"02509021";
		ram_buffer(306) := X"2411FFFF";
		ram_buffer(307) := X"8E650004";
		ram_buffer(308) := X"24060004";
		ram_buffer(309) := X"00052880";
		ram_buffer(310) := X"02052821";
		ram_buffer(311) := X"0C000141";
		ram_buffer(312) := X"00002025";
		ram_buffer(313) := X"8E420000";
		ram_buffer(314) := X"00000000";
		ram_buffer(315) := X"1051FFF7";
		ram_buffer(316) := X"00000000";
		ram_buffer(317) := X"0040F809";
		ram_buffer(318) := X"00000000";
		ram_buffer(319) := X"1000FFE8";
		ram_buffer(320) := X"00000000";
		ram_buffer(321) := X"10C00020";
		ram_buffer(322) := X"00000000";
		ram_buffer(323) := X"27BDFFE0";
		ram_buffer(324) := X"00C53021";
		ram_buffer(325) := X"AFB00010";
		ram_buffer(326) := X"2410FFF0";
		ram_buffer(327) := X"00D01024";
		ram_buffer(328) := X"0046302B";
		ram_buffer(329) := X"AFB20018";
		ram_buffer(330) := X"AFB10014";
		ram_buffer(331) := X"24520010";
		ram_buffer(332) := X"00808825";
		ram_buffer(333) := X"00063100";
		ram_buffer(334) := X"00002025";
		ram_buffer(335) := X"AFBF001C";
		ram_buffer(336) := X"00B08024";
		ram_buffer(337) := X"02469021";
		ram_buffer(338) := X"0C000046";
		ram_buffer(339) := X"2631FF00";
		ram_buffer(340) := X"2403FFF0";
		ram_buffer(341) := X"16500008";
		ram_buffer(342) := X"02032024";
		ram_buffer(343) := X"8FBF001C";
		ram_buffer(344) := X"8FB20018";
		ram_buffer(345) := X"8FB10014";
		ram_buffer(346) := X"8FB00010";
		ram_buffer(347) := X"00402025";
		ram_buffer(348) := X"08000046";
		ram_buffer(349) := X"27BD0020";
		ram_buffer(350) := X"AE240000";
		ram_buffer(351) := X"AC800000";
		ram_buffer(352) := X"1000FFF4";
		ram_buffer(353) := X"26100010";
		ram_buffer(354) := X"03E00008";
		ram_buffer(355) := X"00000000";
		ram_buffer(356) := X"24020001";
		ram_buffer(357) := X"14400002";
		ram_buffer(358) := X"0082001B";
		ram_buffer(359) := X"0007000D";
		ram_buffer(360) := X"00001812";
		ram_buffer(361) := X"0065182B";
		ram_buffer(362) := X"10600006";
		ram_buffer(363) := X"00450018";
		ram_buffer(364) := X"00004025";
		ram_buffer(365) := X"14400006";
		ram_buffer(366) := X"00000000";
		ram_buffer(367) := X"03E00008";
		ram_buffer(368) := X"A0E00000";
		ram_buffer(369) := X"00001012";
		ram_buffer(370) := X"1000FFF2";
		ram_buffer(371) := X"00000000";
		ram_buffer(372) := X"14400002";
		ram_buffer(373) := X"0082001B";
		ram_buffer(374) := X"0007000D";
		ram_buffer(375) := X"00002010";
		ram_buffer(376) := X"00004812";
		ram_buffer(377) := X"00000000";
		ram_buffer(378) := X"00000000";
		ram_buffer(379) := X"14A00002";
		ram_buffer(380) := X"0045001B";
		ram_buffer(381) := X"0007000D";
		ram_buffer(382) := X"00001012";
		ram_buffer(383) := X"15000005";
		ram_buffer(384) := X"292A000A";
		ram_buffer(385) := X"1D200004";
		ram_buffer(386) := X"24EB0001";
		ram_buffer(387) := X"1440FFE9";
		ram_buffer(388) := X"00000000";
		ram_buffer(389) := X"24EB0001";
		ram_buffer(390) := X"15400004";
		ram_buffer(391) := X"24030030";
		ram_buffer(392) := X"14C00002";
		ram_buffer(393) := X"24030037";
		ram_buffer(394) := X"24030057";
		ram_buffer(395) := X"00691821";
		ram_buffer(396) := X"A0E30000";
		ram_buffer(397) := X"25080001";
		ram_buffer(398) := X"1000FFDE";
		ram_buffer(399) := X"01603825";
		ram_buffer(400) := X"27BDFFD8";
		ram_buffer(401) := X"AFB40020";
		ram_buffer(402) := X"AFB3001C";
		ram_buffer(403) := X"AFB20018";
		ram_buffer(404) := X"AFB10014";
		ram_buffer(405) := X"AFBF0024";
		ram_buffer(406) := X"AFB00010";
		ram_buffer(407) := X"00809025";
		ram_buffer(408) := X"00A09825";
		ram_buffer(409) := X"8FB10038";
		ram_buffer(410) := X"10E00002";
		ram_buffer(411) := X"24140020";
		ram_buffer(412) := X"24140030";
		ram_buffer(413) := X"02201025";
		ram_buffer(414) := X"24420001";
		ram_buffer(415) := X"8043FFFF";
		ram_buffer(416) := X"00000000";
		ram_buffer(417) := X"14600009";
		ram_buffer(418) := X"00C08025";
		ram_buffer(419) := X"1A000009";
		ram_buffer(420) := X"02802825";
		ram_buffer(421) := X"0260F809";
		ram_buffer(422) := X"02402025";
		ram_buffer(423) := X"1000FFFB";
		ram_buffer(424) := X"2610FFFF";
		ram_buffer(425) := X"1000FFF4";
		ram_buffer(426) := X"24C6FFFF";
		ram_buffer(427) := X"1CC0FFFD";
		ram_buffer(428) := X"00000000";
		ram_buffer(429) := X"26310001";
		ram_buffer(430) := X"8225FFFF";
		ram_buffer(431) := X"00000000";
		ram_buffer(432) := X"14A00009";
		ram_buffer(433) := X"00000000";
		ram_buffer(434) := X"8FBF0024";
		ram_buffer(435) := X"8FB40020";
		ram_buffer(436) := X"8FB3001C";
		ram_buffer(437) := X"8FB20018";
		ram_buffer(438) := X"8FB10014";
		ram_buffer(439) := X"8FB00010";
		ram_buffer(440) := X"03E00008";
		ram_buffer(441) := X"27BD0028";
		ram_buffer(442) := X"0260F809";
		ram_buffer(443) := X"02402025";
		ram_buffer(444) := X"1000FFF1";
		ram_buffer(445) := X"26310001";
		ram_buffer(446) := X"8C820000";
		ram_buffer(447) := X"00000000";
		ram_buffer(448) := X"24430001";
		ram_buffer(449) := X"AC830000";
		ram_buffer(450) := X"03E00008";
		ram_buffer(451) := X"A0450000";
		ram_buffer(452) := X"27BDFFB8";
		ram_buffer(453) := X"AFB5003C";
		ram_buffer(454) := X"AFB40038";
		ram_buffer(455) := X"AFB30034";
		ram_buffer(456) := X"AFB20030";
		ram_buffer(457) := X"AFB1002C";
		ram_buffer(458) := X"AFB00028";
		ram_buffer(459) := X"AFBF0044";
		ram_buffer(460) := X"AFB60040";
		ram_buffer(461) := X"00809025";
		ram_buffer(462) := X"00A09825";
		ram_buffer(463) := X"00C08825";
		ram_buffer(464) := X"00E08025";
		ram_buffer(465) := X"24140025";
		ram_buffer(466) := X"24150030";
		ram_buffer(467) := X"82250000";
		ram_buffer(468) := X"00000000";
		ram_buffer(469) := X"10A00035";
		ram_buffer(470) := X"00000000";
		ram_buffer(471) := X"10B40006";
		ram_buffer(472) := X"00000000";
		ram_buffer(473) := X"26310001";
		ram_buffer(474) := X"0260F809";
		ram_buffer(475) := X"02402025";
		ram_buffer(476) := X"1000FFF6";
		ram_buffer(477) := X"00000000";
		ram_buffer(478) := X"82260001";
		ram_buffer(479) := X"00000000";
		ram_buffer(480) := X"10D50015";
		ram_buffer(481) := X"240D0001";
		ram_buffer(482) := X"26310002";
		ram_buffer(483) := X"00006825";
		ram_buffer(484) := X"24C2FFD0";
		ram_buffer(485) := X"304200FF";
		ram_buffer(486) := X"2C42000A";
		ram_buffer(487) := X"10400018";
		ram_buffer(488) := X"00006025";
		ram_buffer(489) := X"30C200FF";
		ram_buffer(490) := X"2443FFD0";
		ram_buffer(491) := X"2C63000A";
		ram_buffer(492) := X"1060000C";
		ram_buffer(493) := X"2443FF9F";
		ram_buffer(494) := X"24C3FFD0";
		ram_buffer(495) := X"000C1080";
		ram_buffer(496) := X"004C6021";
		ram_buffer(497) := X"000C6040";
		ram_buffer(498) := X"26310001";
		ram_buffer(499) := X"8226FFFF";
		ram_buffer(500) := X"1000FFF4";
		ram_buffer(501) := X"01836021";
		ram_buffer(502) := X"82260002";
		ram_buffer(503) := X"1000FFEC";
		ram_buffer(504) := X"26310003";
		ram_buffer(505) := X"2C630006";
		ram_buffer(506) := X"1060001A";
		ram_buffer(507) := X"2442FFBF";
		ram_buffer(508) := X"24C3FFA9";
		ram_buffer(509) := X"2862000B";
		ram_buffer(510) := X"1440FFF1";
		ram_buffer(511) := X"000C1080";
		ram_buffer(512) := X"24020063";
		ram_buffer(513) := X"10C20045";
		ram_buffer(514) := X"28C20064";
		ram_buffer(515) := X"10400016";
		ram_buffer(516) := X"24020073";
		ram_buffer(517) := X"10D4004C";
		ram_buffer(518) := X"24020058";
		ram_buffer(519) := X"10C20033";
		ram_buffer(520) := X"00000000";
		ram_buffer(521) := X"14C0FFC9";
		ram_buffer(522) := X"00000000";
		ram_buffer(523) := X"8FBF0044";
		ram_buffer(524) := X"8FB60040";
		ram_buffer(525) := X"8FB5003C";
		ram_buffer(526) := X"8FB40038";
		ram_buffer(527) := X"8FB30034";
		ram_buffer(528) := X"8FB20030";
		ram_buffer(529) := X"8FB1002C";
		ram_buffer(530) := X"8FB00028";
		ram_buffer(531) := X"03E00008";
		ram_buffer(532) := X"27BD0048";
		ram_buffer(533) := X"2C420006";
		ram_buffer(534) := X"1040FFEA";
		ram_buffer(535) := X"24020063";
		ram_buffer(536) := X"1000FFE4";
		ram_buffer(537) := X"24C3FFC9";
		ram_buffer(538) := X"10C20032";
		ram_buffer(539) := X"28C20074";
		ram_buffer(540) := X"10400019";
		ram_buffer(541) := X"24020075";
		ram_buffer(542) := X"24020064";
		ram_buffer(543) := X"14C2FFB3";
		ram_buffer(544) := X"26160004";
		ram_buffer(545) := X"8E040000";
		ram_buffer(546) := X"00000000";
		ram_buffer(547) := X"04810005";
		ram_buffer(548) := X"27A70018";
		ram_buffer(549) := X"2402002D";
		ram_buffer(550) := X"00042023";
		ram_buffer(551) := X"A3A20018";
		ram_buffer(552) := X"27A70019";
		ram_buffer(553) := X"00003025";
		ram_buffer(554) := X"2405000A";
		ram_buffer(555) := X"0C000164";
		ram_buffer(556) := X"00000000";
		ram_buffer(557) := X"27A20018";
		ram_buffer(558) := X"AFA20010";
		ram_buffer(559) := X"01A03825";
		ram_buffer(560) := X"01803025";
		ram_buffer(561) := X"02602825";
		ram_buffer(562) := X"0C000190";
		ram_buffer(563) := X"02402025";
		ram_buffer(564) := X"1000FF9E";
		ram_buffer(565) := X"02C08025";
		ram_buffer(566) := X"10C2000A";
		ram_buffer(567) := X"26160004";
		ram_buffer(568) := X"24020078";
		ram_buffer(569) := X"14C2FF99";
		ram_buffer(570) := X"00000000";
		ram_buffer(571) := X"38C60058";
		ram_buffer(572) := X"26160004";
		ram_buffer(573) := X"27A70018";
		ram_buffer(574) := X"2CC60001";
		ram_buffer(575) := X"10000004";
		ram_buffer(576) := X"24050010";
		ram_buffer(577) := X"27A70018";
		ram_buffer(578) := X"00003025";
		ram_buffer(579) := X"2405000A";
		ram_buffer(580) := X"8E040000";
		ram_buffer(581) := X"1000FFE5";
		ram_buffer(582) := X"00000000";
		ram_buffer(583) := X"82050003";
		ram_buffer(584) := X"02402025";
		ram_buffer(585) := X"0260F809";
		ram_buffer(586) := X"26160004";
		ram_buffer(587) := X"1000FF87";
		ram_buffer(588) := X"02C08025";
		ram_buffer(589) := X"8E020000";
		ram_buffer(590) := X"26160004";
		ram_buffer(591) := X"AFA20010";
		ram_buffer(592) := X"1000FFDF";
		ram_buffer(593) := X"00003825";
		ram_buffer(594) := X"1000FF87";
		ram_buffer(595) := X"24050025";
		ram_buffer(596) := X"AF858014";
		ram_buffer(597) := X"03E00008";
		ram_buffer(598) := X"AF848010";
		ram_buffer(599) := X"27BDFFE0";
		ram_buffer(600) := X"AFA50024";
		ram_buffer(601) := X"AFA60028";
		ram_buffer(602) := X"8F858014";
		ram_buffer(603) := X"00803025";
		ram_buffer(604) := X"8F848010";
		ram_buffer(605) := X"AFA7002C";
		ram_buffer(606) := X"27A70024";
		ram_buffer(607) := X"AFBF001C";
		ram_buffer(608) := X"0C0001C4";
		ram_buffer(609) := X"AFA70010";
		ram_buffer(610) := X"8FBF001C";
		ram_buffer(611) := X"00000000";
		ram_buffer(612) := X"03E00008";
		ram_buffer(613) := X"27BD0020";
		ram_buffer(614) := X"27BDFFE0";
		ram_buffer(615) := X"AFA60028";
		ram_buffer(616) := X"00A03025";
		ram_buffer(617) := X"3C051000";
		ram_buffer(618) := X"AFA40020";
		ram_buffer(619) := X"AFA7002C";
		ram_buffer(620) := X"27A40020";
		ram_buffer(621) := X"27A70028";
		ram_buffer(622) := X"24A506F8";
		ram_buffer(623) := X"AFBF001C";
		ram_buffer(624) := X"0C0001C4";
		ram_buffer(625) := X"AFA70010";
		ram_buffer(626) := X"8FA20020";
		ram_buffer(627) := X"00000000";
		ram_buffer(628) := X"A0400000";
		ram_buffer(629) := X"8FBF001C";
		ram_buffer(630) := X"00000000";
		ram_buffer(631) := X"03E00008";
		ram_buffer(632) := X"27BD0020";
		ram_buffer(633) := X"27BDFFE0";
		ram_buffer(634) := X"AFBF001C";
		ram_buffer(635) := X"AFB10018";
		ram_buffer(636) := X"AFB00014";
		ram_buffer(637) := X"3C031000";
		ram_buffer(638) := X"8C621800";
		ram_buffer(639) := X"3C111000";
		ram_buffer(640) := X"8C420004";
		ram_buffer(641) := X"00608025";
		ram_buffer(642) := X"26311804";
		ram_buffer(643) := X"2C430008";
		ram_buffer(644) := X"14600006";
		ram_buffer(645) := X"00000000";
		ram_buffer(646) := X"8FBF001C";
		ram_buffer(647) := X"8FB10018";
		ram_buffer(648) := X"8FB00014";
		ram_buffer(649) := X"03E00008";
		ram_buffer(650) := X"27BD0020";
		ram_buffer(651) := X"000210C0";
		ram_buffer(652) := X"02221021";
		ram_buffer(653) := X"8C430000";
		ram_buffer(654) := X"8C440004";
		ram_buffer(655) := X"0060F809";
		ram_buffer(656) := X"00000000";
		ram_buffer(657) := X"8E021800";
		ram_buffer(658) := X"00000000";
		ram_buffer(659) := X"8C420004";
		ram_buffer(660) := X"1000FFEF";
		ram_buffer(661) := X"2C430008";
		ram_buffer(662) := X"8F828024";
		ram_buffer(663) := X"00000000";
		ram_buffer(664) := X"8C440004";
		ram_buffer(665) := X"8F82801C";
		ram_buffer(666) := X"8F838018";
		ram_buffer(667) := X"24420001";
		ram_buffer(668) := X"304201FF";
		ram_buffer(669) := X"10430008";
		ram_buffer(670) := X"00000000";
		ram_buffer(671) := X"8F83801C";
		ram_buffer(672) := X"3C051000";
		ram_buffer(673) := X"24A51600";
		ram_buffer(674) := X"308400FF";
		ram_buffer(675) := X"00651821";
		ram_buffer(676) := X"A0640000";
		ram_buffer(677) := X"AF82801C";
		ram_buffer(678) := X"03E00008";
		ram_buffer(679) := X"00000000";
		ram_buffer(680) := X"8F838024";
		ram_buffer(681) := X"00000000";
		ram_buffer(682) := X"8C620000";
		ram_buffer(683) := X"00000000";
		ram_buffer(684) := X"30420002";
		ram_buffer(685) := X"1040FFFC";
		ram_buffer(686) := X"00000000";
		ram_buffer(687) := X"AC650008";
		ram_buffer(688) := X"03E00008";
		ram_buffer(689) := X"00000000";
		ram_buffer(690) := X"3C022000";
		ram_buffer(691) := X"AF828028";
		ram_buffer(692) := X"3C022004";
		ram_buffer(693) := X"AF828024";
		ram_buffer(694) := X"3C022003";
		ram_buffer(695) := X"AF828020";
		ram_buffer(696) := X"3C031000";
		ram_buffer(697) := X"3C022001";
		ram_buffer(698) := X"27BDFFE8";
		ram_buffer(699) := X"AC621800";
		ram_buffer(700) := X"3C041000";
		ram_buffer(701) := X"3C021000";
		ram_buffer(702) := X"24421804";
		ram_buffer(703) := X"AFBF0014";
		ram_buffer(704) := X"AFB00010";
		ram_buffer(705) := X"24841844";
		ram_buffer(706) := X"24420008";
		ram_buffer(707) := X"1444FFFE";
		ram_buffer(708) := X"AC40FFF8";
		ram_buffer(709) := X"3C021000";
		ram_buffer(710) := X"24701800";
		ram_buffer(711) := X"24420A58";
		ram_buffer(712) := X"AE020014";
		ram_buffer(713) := X"AE000018";
		ram_buffer(714) := X"3C06F000";
		ram_buffer(715) := X"8CC40004";
		ram_buffer(716) := X"3C051000";
		ram_buffer(717) := X"00041100";
		ram_buffer(718) := X"00441021";
		ram_buffer(719) := X"00021080";
		ram_buffer(720) := X"3C041000";
		ram_buffer(721) := X"24840EE0";
		ram_buffer(722) := X"24420004";
		ram_buffer(723) := X"00821021";
		ram_buffer(724) := X"24A509E4";
		ram_buffer(725) := X"AC450008";
		ram_buffer(726) := X"AC40000C";
		ram_buffer(727) := X"8C631800";
		ram_buffer(728) := X"00000000";
		ram_buffer(729) := X"8C620000";
		ram_buffer(730) := X"00000000";
		ram_buffer(731) := X"34420004";
		ram_buffer(732) := X"AC620000";
		ram_buffer(733) := X"8CC30004";
		ram_buffer(734) := X"00000000";
		ram_buffer(735) := X"00031100";
		ram_buffer(736) := X"00431021";
		ram_buffer(737) := X"00021080";
		ram_buffer(738) := X"00441021";
		ram_buffer(739) := X"8C430000";
		ram_buffer(740) := X"24060004";
		ram_buffer(741) := X"8C620000";
		ram_buffer(742) := X"27858028";
		ram_buffer(743) := X"34420002";
		ram_buffer(744) := X"AC620000";
		ram_buffer(745) := X"0C000141";
		ram_buffer(746) := X"24040004";
		ram_buffer(747) := X"24060004";
		ram_buffer(748) := X"27858024";
		ram_buffer(749) := X"0C000141";
		ram_buffer(750) := X"24040004";
		ram_buffer(751) := X"24060004";
		ram_buffer(752) := X"27858020";
		ram_buffer(753) := X"0C000141";
		ram_buffer(754) := X"24040004";
		ram_buffer(755) := X"24060044";
		ram_buffer(756) := X"02002825";
		ram_buffer(757) := X"0C000141";
		ram_buffer(758) := X"24040004";
		ram_buffer(759) := X"3C021000";
		ram_buffer(760) := X"2442003C";
		ram_buffer(761) := X"2403003C";
		ram_buffer(762) := X"10430007";
		ram_buffer(763) := X"00000000";
		ram_buffer(764) := X"0C000049";
		ram_buffer(765) := X"00000000";
		ram_buffer(766) := X"24060010";
		ram_buffer(767) := X"2405003C";
		ram_buffer(768) := X"0C000141";
		ram_buffer(769) := X"24040004";
		ram_buffer(770) := X"8FBF0014";
		ram_buffer(771) := X"8FB00010";
		ram_buffer(772) := X"24040001";
		ram_buffer(773) := X"08000046";
		ram_buffer(774) := X"27BD0018";
		ram_buffer(775) := X"27BDFFE8";
		ram_buffer(776) := X"24060004";
		ram_buffer(777) := X"27858028";
		ram_buffer(778) := X"AFBF0014";
		ram_buffer(779) := X"0C000141";
		ram_buffer(780) := X"00002025";
		ram_buffer(781) := X"24060004";
		ram_buffer(782) := X"27858024";
		ram_buffer(783) := X"0C000141";
		ram_buffer(784) := X"00002025";
		ram_buffer(785) := X"24060004";
		ram_buffer(786) := X"27858020";
		ram_buffer(787) := X"0C000141";
		ram_buffer(788) := X"00002025";
		ram_buffer(789) := X"3C051000";
		ram_buffer(790) := X"24060044";
		ram_buffer(791) := X"24A51800";
		ram_buffer(792) := X"0C000141";
		ram_buffer(793) := X"00002025";
		ram_buffer(794) := X"3C051000";
		ram_buffer(795) := X"24A50AA0";
		ram_buffer(796) := X"0C000254";
		ram_buffer(797) := X"00002025";
		ram_buffer(798) := X"3C021000";
		ram_buffer(799) := X"2442003C";
		ram_buffer(800) := X"2403003C";
		ram_buffer(801) := X"10430004";
		ram_buffer(802) := X"24060010";
		ram_buffer(803) := X"2405003C";
		ram_buffer(804) := X"0C000141";
		ram_buffer(805) := X"00002025";
		ram_buffer(806) := X"8FBF0014";
		ram_buffer(807) := X"24040001";
		ram_buffer(808) := X"08000046";
		ram_buffer(809) := X"27BD0018";
		ram_buffer(810) := X"27BDFFE8";
		ram_buffer(811) := X"AFBF0014";
		ram_buffer(812) := X"0C000046";
		ram_buffer(813) := X"00002025";
		ram_buffer(814) := X"3C021000";
		ram_buffer(815) := X"8C431800";
		ram_buffer(816) := X"2404FFFB";
		ram_buffer(817) := X"8C620000";
		ram_buffer(818) := X"00000000";
		ram_buffer(819) := X"00441024";
		ram_buffer(820) := X"AC620000";
		ram_buffer(821) := X"3C02F000";
		ram_buffer(822) := X"8C430004";
		ram_buffer(823) := X"00000000";
		ram_buffer(824) := X"00031100";
		ram_buffer(825) := X"00431021";
		ram_buffer(826) := X"3C031000";
		ram_buffer(827) := X"24630EE0";
		ram_buffer(828) := X"00021080";
		ram_buffer(829) := X"00431021";
		ram_buffer(830) := X"8C430000";
		ram_buffer(831) := X"8FBF0014";
		ram_buffer(832) := X"8C620000";
		ram_buffer(833) := X"2404FFFD";
		ram_buffer(834) := X"00441024";
		ram_buffer(835) := X"AC620000";
		ram_buffer(836) := X"03E00008";
		ram_buffer(837) := X"27BD0018";
		ram_buffer(838) := X"8F838024";
		ram_buffer(839) := X"00000000";
		ram_buffer(840) := X"8C620000";
		ram_buffer(841) := X"00000000";
		ram_buffer(842) := X"30420002";
		ram_buffer(843) := X"1040FFFC";
		ram_buffer(844) := X"00000000";
		ram_buffer(845) := X"AC640008";
		ram_buffer(846) := X"03E00008";
		ram_buffer(847) := X"00000000";
		ram_buffer(848) := X"27BDFFE8";
		ram_buffer(849) := X"AFBF0014";
		ram_buffer(850) := X"AFB00010";
		ram_buffer(851) := X"0C000046";
		ram_buffer(852) := X"00002025";
		ram_buffer(853) := X"8F83801C";
		ram_buffer(854) := X"8F828018";
		ram_buffer(855) := X"00000000";
		ram_buffer(856) := X"14620005";
		ram_buffer(857) := X"00000000";
		ram_buffer(858) := X"0C000046";
		ram_buffer(859) := X"24040001";
		ram_buffer(860) := X"1000FFF6";
		ram_buffer(861) := X"00000000";
		ram_buffer(862) := X"8F828018";
		ram_buffer(863) := X"3C031000";
		ram_buffer(864) := X"24631600";
		ram_buffer(865) := X"00431021";
		ram_buffer(866) := X"90500000";
		ram_buffer(867) := X"8F828018";
		ram_buffer(868) := X"24040001";
		ram_buffer(869) := X"24420001";
		ram_buffer(870) := X"304201FF";
		ram_buffer(871) := X"AF828018";
		ram_buffer(872) := X"0C000046";
		ram_buffer(873) := X"321000FF";
		ram_buffer(874) := X"8FBF0014";
		ram_buffer(875) := X"02001025";
		ram_buffer(876) := X"8FB00010";
		ram_buffer(877) := X"03E00008";
		ram_buffer(878) := X"27BD0018";
		ram_buffer(879) := X"27BDFFE8";
		ram_buffer(880) := X"00803025";
		ram_buffer(881) := X"24050004";
		ram_buffer(882) := X"AFBF0014";
		ram_buffer(883) := X"0C000346";
		ram_buffer(884) := X"30C400FF";
		ram_buffer(885) := X"24A5FFFF";
		ram_buffer(886) := X"14A0FFFC";
		ram_buffer(887) := X"00063202";
		ram_buffer(888) := X"8FBF0014";
		ram_buffer(889) := X"00000000";
		ram_buffer(890) := X"03E00008";
		ram_buffer(891) := X"27BD0018";
		ram_buffer(892) := X"27BDFFE0";
		ram_buffer(893) := X"AFB20018";
		ram_buffer(894) := X"AFB10014";
		ram_buffer(895) := X"AFB00010";
		ram_buffer(896) := X"AFBF001C";
		ram_buffer(897) := X"00008025";
		ram_buffer(898) := X"00008825";
		ram_buffer(899) := X"24120020";
		ram_buffer(900) := X"0C000350";
		ram_buffer(901) := X"00000000";
		ram_buffer(902) := X"02021004";
		ram_buffer(903) := X"26100008";
		ram_buffer(904) := X"1612FFFB";
		ram_buffer(905) := X"02228825";
		ram_buffer(906) := X"8FBF001C";
		ram_buffer(907) := X"02201025";
		ram_buffer(908) := X"8FB20018";
		ram_buffer(909) := X"8FB10014";
		ram_buffer(910) := X"8FB00010";
		ram_buffer(911) := X"03E00008";
		ram_buffer(912) := X"27BD0020";
		ram_buffer(913) := X"8F828020";
		ram_buffer(914) := X"00000000";
		ram_buffer(915) := X"03E00008";
		ram_buffer(916) := X"AC440008";
		ram_buffer(917) := X"3C04F000";
		ram_buffer(918) := X"8C820004";
		ram_buffer(919) := X"00000000";
		ram_buffer(920) := X"24420001";
		ram_buffer(921) := X"8F838028";
		ram_buffer(922) := X"00000000";
		ram_buffer(923) := X"AC620000";
		ram_buffer(924) := X"8F838028";
		ram_buffer(925) := X"00000000";
		ram_buffer(926) := X"8C630000";
		ram_buffer(927) := X"00000000";
		ram_buffer(928) := X"1443FFF5";
		ram_buffer(929) := X"00000000";
		ram_buffer(930) := X"03E00008";
		ram_buffer(931) := X"00000000";
		ram_buffer(932) := X"8F838028";
		ram_buffer(933) := X"3C02F000";
		ram_buffer(934) := X"8C420004";
		ram_buffer(935) := X"00000000";
		ram_buffer(936) := X"24420001";
		ram_buffer(937) := X"03E00008";
		ram_buffer(938) := X"AC620000";
		ram_buffer(939) := X"00000000";
		ram_buffer(940) := X"00000100";
		ram_buffer(941) := X"01010001";
		ram_buffer(942) := X"00000000";
		ram_buffer(943) := X"00000000";
		ram_buffer(944) := X"00000000";
		ram_buffer(945) := X"00000000";
		ram_buffer(946) := X"FFFFFFFF";
		ram_buffer(947) := X"FFFFFFFF";
		ram_buffer(948) := X"FFFFFFFF";
		ram_buffer(949) := X"FFFFFFFF";
		ram_buffer(950) := X"FFFFFFFF";
		ram_buffer(951) := X"FFFFFFFF";
		ram_buffer(952) := X"FFFFFFFF";
		ram_buffer(953) := X"00000000";
		ram_buffer(954) := X"00000000";
		ram_buffer(955) := X"00000000";
		ram_buffer(956) := X"00000000";
		ram_buffer(957) := X"00000000";
		ram_buffer(958) := X"00000000";
		ram_buffer(959) := X"00000000";
		ram_buffer(960) := X"00000000";
		ram_buffer(961) := X"00000000";
		ram_buffer(962) := X"00000000";
		ram_buffer(963) := X"00000000";
		ram_buffer(964) := X"00000000";
		ram_buffer(965) := X"00000000";
		ram_buffer(966) := X"00000000";
		ram_buffer(967) := X"00000000";
		ram_buffer(968) := X"00000000";
		ram_buffer(969) := X"FFFFFFFF";
		ram_buffer(970) := X"00000000";
		ram_buffer(971) := X"00000000";
		ram_buffer(972) := X"00000000";
		ram_buffer(973) := X"00000000";
		ram_buffer(974) := X"00000000";
		ram_buffer(975) := X"00000000";
		ram_buffer(976) := X"00000000";
		ram_buffer(977) := X"00000000";
		ram_buffer(978) := X"00000000";
		ram_buffer(979) := X"00000000";
		ram_buffer(980) := X"00000000";
		ram_buffer(981) := X"00000000";
		ram_buffer(982) := X"00000000";
		ram_buffer(983) := X"00000000";
		ram_buffer(984) := X"00000000";
		ram_buffer(985) := X"00000000";
		ram_buffer(986) := X"FFFFFFFF";
		ram_buffer(987) := X"00000000";
		ram_buffer(988) := X"00000000";
		ram_buffer(989) := X"00000000";
		ram_buffer(990) := X"00000000";
		ram_buffer(991) := X"00000000";
		ram_buffer(992) := X"00000000";
		ram_buffer(993) := X"00000000";
		ram_buffer(994) := X"00000000";
		ram_buffer(995) := X"00000000";
		ram_buffer(996) := X"00000000";
		ram_buffer(997) := X"00000000";
		ram_buffer(998) := X"00000000";
		ram_buffer(999) := X"00000000";
		ram_buffer(1000) := X"00000000";
		ram_buffer(1001) := X"00000000";
		ram_buffer(1002) := X"00000000";
		return ram_buffer;
	end;
end;
