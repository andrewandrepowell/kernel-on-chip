
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

package nexys4_pack is

    constant data_out_width : integer := 16;
    constant data_in_width : integer := 16;

end package;