library ieee;
use ieee.std_logic_1164.all;

package main_pack is

	constant cpu_width : integer := 32;
	constant ram_size : integer := 306;
	subtype word_type is std_logic_vector(cpu_width-1 downto 0);
	type ram_type is array(0 to ram_size-1) of word_type;
	function load_hex return ram_type;

end package;

package body main_pack is

	function load_hex return ram_type is
		variable ram_buffer : ram_type := (others=>(others=>'0'));
	begin
		ram_buffer(0) := X"3C1C1001";
		ram_buffer(1) := X"279C84C0";
		ram_buffer(2) := X"3C1D1000";
		ram_buffer(3) := X"27BD04E8";
		ram_buffer(4) := X"0C00009F";
		ram_buffer(5) := X"00000000";
		ram_buffer(6) := X"23BDFF98";
		ram_buffer(7) := X"AFA10010";
		ram_buffer(8) := X"AFA20014";
		ram_buffer(9) := X"AFA30018";
		ram_buffer(10) := X"AFA4001C";
		ram_buffer(11) := X"AFA50020";
		ram_buffer(12) := X"AFA60024";
		ram_buffer(13) := X"AFA70028";
		ram_buffer(14) := X"AFA8002C";
		ram_buffer(15) := X"AFA90030";
		ram_buffer(16) := X"AFAA0034";
		ram_buffer(17) := X"AFAB0038";
		ram_buffer(18) := X"AFAC003C";
		ram_buffer(19) := X"AFAD0040";
		ram_buffer(20) := X"AFAE0044";
		ram_buffer(21) := X"AFAF0048";
		ram_buffer(22) := X"AFB8004C";
		ram_buffer(23) := X"AFB90050";
		ram_buffer(24) := X"AFBF0054";
		ram_buffer(25) := X"0C000079";
		ram_buffer(26) := X"23A50000";
		ram_buffer(27) := X"8FA10010";
		ram_buffer(28) := X"8FA20014";
		ram_buffer(29) := X"8FA30018";
		ram_buffer(30) := X"8FA4001C";
		ram_buffer(31) := X"8FA50020";
		ram_buffer(32) := X"8FA60024";
		ram_buffer(33) := X"8FA70028";
		ram_buffer(34) := X"8FA8002C";
		ram_buffer(35) := X"8FA90030";
		ram_buffer(36) := X"8FAA0034";
		ram_buffer(37) := X"8FAB0038";
		ram_buffer(38) := X"8FAC003C";
		ram_buffer(39) := X"8FAD0040";
		ram_buffer(40) := X"8FAE0044";
		ram_buffer(41) := X"8FAF0048";
		ram_buffer(42) := X"8FB8004C";
		ram_buffer(43) := X"8FB90050";
		ram_buffer(44) := X"8FBF0054";
		ram_buffer(45) := X"8FBA0058";
		ram_buffer(46) := X"8FBB005C";
		ram_buffer(47) := X"03600011";
		ram_buffer(48) := X"8FBB0060";
		ram_buffer(49) := X"03600013";
		ram_buffer(50) := X"23BD0068";
		ram_buffer(51) := X"341B0001";
		ram_buffer(52) := X"03400008";
		ram_buffer(53) := X"409B6000";
		ram_buffer(54) := X"40026000";
		ram_buffer(55) := X"03E00008";
		ram_buffer(56) := X"40846000";
		ram_buffer(57) := X"3C051000";
		ram_buffer(58) := X"24A50110";
		ram_buffer(59) := X"8CA60000";
		ram_buffer(60) := X"AC06003C";
		ram_buffer(61) := X"8CA60004";
		ram_buffer(62) := X"AC060040";
		ram_buffer(63) := X"8CA60008";
		ram_buffer(64) := X"AC060044";
		ram_buffer(65) := X"8CA6000C";
		ram_buffer(66) := X"03E00008";
		ram_buffer(67) := X"AC060048";
		ram_buffer(68) := X"3C1A1000";
		ram_buffer(69) := X"375A0018";
		ram_buffer(70) := X"03400008";
		ram_buffer(71) := X"00000000";
		ram_buffer(72) := X"00850019";
		ram_buffer(73) := X"00001012";
		ram_buffer(74) := X"00002010";
		ram_buffer(75) := X"03E00008";
		ram_buffer(76) := X"ACC40000";
		ram_buffer(77) := X"0000000C";
		ram_buffer(78) := X"03E00008";
		ram_buffer(79) := X"00000000";
		ram_buffer(80) := X"AC900000";
		ram_buffer(81) := X"AC910004";
		ram_buffer(82) := X"AC920008";
		ram_buffer(83) := X"AC93000C";
		ram_buffer(84) := X"AC940010";
		ram_buffer(85) := X"AC950014";
		ram_buffer(86) := X"AC960018";
		ram_buffer(87) := X"AC97001C";
		ram_buffer(88) := X"AC9E0020";
		ram_buffer(89) := X"AC9C0024";
		ram_buffer(90) := X"AC9D0028";
		ram_buffer(91) := X"AC9F002C";
		ram_buffer(92) := X"03E00008";
		ram_buffer(93) := X"34020000";
		ram_buffer(94) := X"8C900000";
		ram_buffer(95) := X"8C910004";
		ram_buffer(96) := X"8C920008";
		ram_buffer(97) := X"8C93000C";
		ram_buffer(98) := X"8C940010";
		ram_buffer(99) := X"8C950014";
		ram_buffer(100) := X"8C960018";
		ram_buffer(101) := X"8C97001C";
		ram_buffer(102) := X"8C9E0020";
		ram_buffer(103) := X"8C9C0024";
		ram_buffer(104) := X"8C9D0028";
		ram_buffer(105) := X"8C9F002C";
		ram_buffer(106) := X"03E00008";
		ram_buffer(107) := X"34A20000";
		ram_buffer(108) := X"1000FFFF";
		ram_buffer(109) := X"00000000";
		ram_buffer(110) := X"3C02F000";
		ram_buffer(111) := X"8C420004";
		ram_buffer(112) := X"3C031000";
		ram_buffer(113) := X"246303F0";
		ram_buffer(114) := X"00021080";
		ram_buffer(115) := X"00431021";
		ram_buffer(116) := X"8C420000";
		ram_buffer(117) := X"24030002";
		ram_buffer(118) := X"AC430000";
		ram_buffer(119) := X"03E00008";
		ram_buffer(120) := X"00000000";
		ram_buffer(121) := X"3C02F000";
		ram_buffer(122) := X"8C430004";
		ram_buffer(123) := X"27BDFFE0";
		ram_buffer(124) := X"00031100";
		ram_buffer(125) := X"00431021";
		ram_buffer(126) := X"AFB10014";
		ram_buffer(127) := X"3C111000";
		ram_buffer(128) := X"00021080";
		ram_buffer(129) := X"263103FC";
		ram_buffer(130) := X"AFB20018";
		ram_buffer(131) := X"24520004";
		ram_buffer(132) := X"02221021";
		ram_buffer(133) := X"8C430000";
		ram_buffer(134) := X"AFB00010";
		ram_buffer(135) := X"8C630004";
		ram_buffer(136) := X"AFBF001C";
		ram_buffer(137) := X"00408025";
		ram_buffer(138) := X"2C620008";
		ram_buffer(139) := X"14400007";
		ram_buffer(140) := X"00000000";
		ram_buffer(141) := X"8FBF001C";
		ram_buffer(142) := X"8FB20018";
		ram_buffer(143) := X"8FB10014";
		ram_buffer(144) := X"8FB00010";
		ram_buffer(145) := X"03E00008";
		ram_buffer(146) := X"27BD0020";
		ram_buffer(147) := X"000318C0";
		ram_buffer(148) := X"00721821";
		ram_buffer(149) := X"02231821";
		ram_buffer(150) := X"8C620000";
		ram_buffer(151) := X"8C640004";
		ram_buffer(152) := X"0040F809";
		ram_buffer(153) := X"00000000";
		ram_buffer(154) := X"8E020000";
		ram_buffer(155) := X"00000000";
		ram_buffer(156) := X"8C430004";
		ram_buffer(157) := X"1000FFED";
		ram_buffer(158) := X"2C620008";
		ram_buffer(159) := X"3C05F000";
		ram_buffer(160) := X"8CA20004";
		ram_buffer(161) := X"27BDFFE8";
		ram_buffer(162) := X"00021240";
		ram_buffer(163) := X"244301E8";
		ram_buffer(164) := X"3C021000";
		ram_buffer(165) := X"24420544";
		ram_buffer(166) := X"00431021";
		ram_buffer(167) := X"AFBF0014";
		ram_buffer(168) := X"0040E825";
		ram_buffer(169) := X"8CA70004";
		ram_buffer(170) := X"8CA20004";
		ram_buffer(171) := X"3C031000";
		ram_buffer(172) := X"246303F0";
		ram_buffer(173) := X"00021080";
		ram_buffer(174) := X"00431021";
		ram_buffer(175) := X"00072100";
		ram_buffer(176) := X"3C03F002";
		ram_buffer(177) := X"AC430000";
		ram_buffer(178) := X"00871021";
		ram_buffer(179) := X"3C031000";
		ram_buffer(180) := X"00021080";
		ram_buffer(181) := X"246303FC";
		ram_buffer(182) := X"00432821";
		ram_buffer(183) := X"24420004";
		ram_buffer(184) := X"3C06F001";
		ram_buffer(185) := X"00621021";
		ram_buffer(186) := X"ACA60000";
		ram_buffer(187) := X"24A60044";
		ram_buffer(188) := X"00402825";
		ram_buffer(189) := X"14C50021";
		ram_buffer(190) := X"24A50008";
		ram_buffer(191) := X"3C051000";
		ram_buffer(192) := X"24A501B8";
		ram_buffer(193) := X"AC450000";
		ram_buffer(194) := X"AC400004";
		ram_buffer(195) := X"00872021";
		ram_buffer(196) := X"00042080";
		ram_buffer(197) := X"00641821";
		ram_buffer(198) := X"8C620000";
		ram_buffer(199) := X"24030001";
		ram_buffer(200) := X"0C000039";
		ram_buffer(201) := X"AC430000";
		ram_buffer(202) := X"3C02F000";
		ram_buffer(203) := X"8C420004";
		ram_buffer(204) := X"00000000";
		ram_buffer(205) := X"1440000D";
		ram_buffer(206) := X"27868008";
		ram_buffer(207) := X"27828684";
		ram_buffer(208) := X"14C20010";
		ram_buffer(209) := X"24C60004";
		ram_buffer(210) := X"24C6FFFC";
		ram_buffer(211) := X"27828008";
		ram_buffer(212) := X"24C60004";
		ram_buffer(213) := X"00C23023";
		ram_buffer(214) := X"00402825";
		ram_buffer(215) := X"0C0000E3";
		ram_buffer(216) := X"24040004";
		ram_buffer(217) := X"0C00006C";
		ram_buffer(218) := X"00000000";
		ram_buffer(219) := X"0C000036";
		ram_buffer(220) := X"24040001";
		ram_buffer(221) := X"1000FFFF";
		ram_buffer(222) := X"00000000";
		ram_buffer(223) := X"1000FFDD";
		ram_buffer(224) := X"ACA0FFF8";
		ram_buffer(225) := X"1000FFEE";
		ram_buffer(226) := X"ACC0FFFC";
		ram_buffer(227) := X"10C0000C";
		ram_buffer(228) := X"00C53021";
		ram_buffer(229) := X"2402FFF0";
		ram_buffer(230) := X"00C21824";
		ram_buffer(231) := X"0066302B";
		ram_buffer(232) := X"00A22824";
		ram_buffer(233) := X"00063100";
		ram_buffer(234) := X"24620010";
		ram_buffer(235) := X"00463021";
		ram_buffer(236) := X"2484FF00";
		ram_buffer(237) := X"2402FFF0";
		ram_buffer(238) := X"14C50003";
		ram_buffer(239) := X"00A21824";
		ram_buffer(240) := X"03E00008";
		ram_buffer(241) := X"00000000";
		ram_buffer(242) := X"AC830000";
		ram_buffer(243) := X"AC600000";
		ram_buffer(244) := X"1000FFF9";
		ram_buffer(245) := X"24A50010";
		ram_buffer(246) := X"00000100";
		ram_buffer(247) := X"01010001";
		ram_buffer(248) := X"00000000";
		ram_buffer(249) := X"00000000";
		ram_buffer(250) := X"00000000";
		ram_buffer(251) := X"00000000";
		ram_buffer(252) := X"FFFFFFFF";
		ram_buffer(253) := X"FFFFFFFF";
		ram_buffer(254) := X"FFFFFFFF";
		ram_buffer(255) := X"FFFFFFFF";
		ram_buffer(256) := X"00000000";
		ram_buffer(257) := X"00000000";
		ram_buffer(258) := X"00000000";
		ram_buffer(259) := X"00000000";
		ram_buffer(260) := X"00000000";
		ram_buffer(261) := X"00000000";
		ram_buffer(262) := X"00000000";
		ram_buffer(263) := X"00000000";
		ram_buffer(264) := X"00000000";
		ram_buffer(265) := X"00000000";
		ram_buffer(266) := X"00000000";
		ram_buffer(267) := X"00000000";
		ram_buffer(268) := X"00000000";
		ram_buffer(269) := X"00000000";
		ram_buffer(270) := X"00000000";
		ram_buffer(271) := X"00000000";
		ram_buffer(272) := X"FFFFFFFF";
		ram_buffer(273) := X"00000000";
		ram_buffer(274) := X"00000000";
		ram_buffer(275) := X"00000000";
		ram_buffer(276) := X"00000000";
		ram_buffer(277) := X"00000000";
		ram_buffer(278) := X"00000000";
		ram_buffer(279) := X"00000000";
		ram_buffer(280) := X"00000000";
		ram_buffer(281) := X"00000000";
		ram_buffer(282) := X"00000000";
		ram_buffer(283) := X"00000000";
		ram_buffer(284) := X"00000000";
		ram_buffer(285) := X"00000000";
		ram_buffer(286) := X"00000000";
		ram_buffer(287) := X"00000000";
		ram_buffer(288) := X"00000000";
		ram_buffer(289) := X"FFFFFFFF";
		ram_buffer(290) := X"00000000";
		ram_buffer(291) := X"00000000";
		ram_buffer(292) := X"00000000";
		ram_buffer(293) := X"00000000";
		ram_buffer(294) := X"00000000";
		ram_buffer(295) := X"00000000";
		ram_buffer(296) := X"00000000";
		ram_buffer(297) := X"00000000";
		ram_buffer(298) := X"00000000";
		ram_buffer(299) := X"00000000";
		ram_buffer(300) := X"00000000";
		ram_buffer(301) := X"00000000";
		ram_buffer(302) := X"00000000";
		ram_buffer(303) := X"00000000";
		ram_buffer(304) := X"00000000";
		ram_buffer(305) := X"00000000";
		return ram_buffer;
	end;
end;
